magic
tech sky130A
magscale 1 2
timestamp 1654035601
<< viali >>
rect 1409 57409 1443 57443
rect 10609 57409 10643 57443
rect 33793 57409 33827 57443
rect 57161 57409 57195 57443
rect 1685 57341 1719 57375
rect 10425 57273 10459 57307
rect 2881 57205 2915 57239
rect 4077 57205 4111 57239
rect 17969 57205 18003 57239
rect 31493 57205 31527 57239
rect 32321 57205 32355 57239
rect 33609 57205 33643 57239
rect 35909 57205 35943 57239
rect 56057 57205 56091 57239
rect 56701 57205 56735 57239
rect 57253 57205 57287 57239
rect 58081 57205 58115 57239
rect 3801 56865 3835 56899
rect 4261 56865 4295 56899
rect 56333 56865 56367 56899
rect 57989 56865 58023 56899
rect 2237 56797 2271 56831
rect 2881 56797 2915 56831
rect 6469 56797 6503 56831
rect 7665 56797 7699 56831
rect 13461 56797 13495 56831
rect 16037 56797 16071 56831
rect 17417 56797 17451 56831
rect 18245 56797 18279 56831
rect 22569 56797 22603 56831
rect 27261 56797 27295 56831
rect 27905 56797 27939 56831
rect 28365 56797 28399 56831
rect 30205 56797 30239 56831
rect 30665 56797 30699 56831
rect 31309 56797 31343 56831
rect 35633 56797 35667 56831
rect 40049 56797 40083 56831
rect 42257 56797 42291 56831
rect 42901 56797 42935 56831
rect 46489 56797 46523 56831
rect 50353 56797 50387 56831
rect 55873 56797 55907 56831
rect 3985 56729 4019 56763
rect 30757 56729 30791 56763
rect 31493 56729 31527 56763
rect 33149 56729 33183 56763
rect 35817 56729 35851 56763
rect 37473 56729 37507 56763
rect 56517 56729 56551 56763
rect 17509 56661 17543 56695
rect 22385 56661 22419 56695
rect 27077 56661 27111 56695
rect 28457 56661 28491 56695
rect 4353 56457 4387 56491
rect 22201 56457 22235 56491
rect 24409 56457 24443 56491
rect 27353 56457 27387 56491
rect 23274 56389 23308 56423
rect 28181 56389 28215 56423
rect 44465 56389 44499 56423
rect 55689 56389 55723 56423
rect 57989 56389 58023 56423
rect 1961 56321 1995 56355
rect 4261 56321 4295 56355
rect 6377 56321 6411 56355
rect 8677 56321 8711 56355
rect 13277 56321 13311 56355
rect 16773 56321 16807 56355
rect 22017 56321 22051 56355
rect 26249 56321 26283 56355
rect 27169 56321 27203 56355
rect 27997 56321 28031 56355
rect 30849 56321 30883 56355
rect 32137 56321 32171 56355
rect 39681 56321 39715 56355
rect 42625 56321 42659 56355
rect 46673 56321 46707 56355
rect 49525 56321 49559 56355
rect 55505 56321 55539 56355
rect 57897 56321 57931 56355
rect 2145 56253 2179 56287
rect 2789 56253 2823 56287
rect 6561 56253 6595 56287
rect 7021 56253 7055 56287
rect 8861 56253 8895 56287
rect 9137 56253 9171 56287
rect 13461 56253 13495 56287
rect 13829 56253 13863 56287
rect 16957 56253 16991 56287
rect 17417 56253 17451 56287
rect 19073 56253 19107 56287
rect 19257 56253 19291 56287
rect 19533 56253 19567 56287
rect 21833 56253 21867 56287
rect 23029 56253 23063 56287
rect 26065 56253 26099 56287
rect 26985 56253 27019 56287
rect 28457 56253 28491 56287
rect 32321 56253 32355 56287
rect 32873 56253 32907 56287
rect 39865 56253 39899 56287
rect 40601 56253 40635 56287
rect 42809 56253 42843 56287
rect 49709 56253 49743 56287
rect 50353 56253 50387 56287
rect 56701 56253 56735 56287
rect 26433 56117 26467 56151
rect 30941 56117 30975 56151
rect 36001 56117 36035 56151
rect 46765 56117 46799 56151
rect 7481 55913 7515 55947
rect 9045 55913 9079 55947
rect 13093 55913 13127 55947
rect 50261 55913 50295 55947
rect 19441 55845 19475 55879
rect 20453 55845 20487 55879
rect 32413 55845 32447 55879
rect 35173 55845 35207 55879
rect 40141 55845 40175 55879
rect 15761 55777 15795 55811
rect 16221 55777 16255 55811
rect 24961 55777 24995 55811
rect 30021 55777 30055 55811
rect 30481 55777 30515 55811
rect 42441 55777 42475 55811
rect 43821 55777 43855 55811
rect 46213 55777 46247 55811
rect 46397 55777 46431 55811
rect 47041 55777 47075 55811
rect 54769 55777 54803 55811
rect 56333 55777 56367 55811
rect 56793 55777 56827 55811
rect 1501 55709 1535 55743
rect 2605 55709 2639 55743
rect 3801 55709 3835 55743
rect 7389 55709 7423 55743
rect 8953 55709 8987 55743
rect 13001 55709 13035 55743
rect 15117 55709 15151 55743
rect 20913 55709 20947 55743
rect 21005 55709 21039 55743
rect 21833 55709 21867 55743
rect 21925 55709 21959 55743
rect 22753 55709 22787 55743
rect 27077 55709 27111 55743
rect 27333 55709 27367 55743
rect 32321 55709 32355 55743
rect 33149 55709 33183 55743
rect 35081 55709 35115 55743
rect 35725 55709 35759 55743
rect 40049 55709 40083 55743
rect 50169 55709 50203 55743
rect 52929 55709 52963 55743
rect 55689 55709 55723 55743
rect 2053 55641 2087 55675
rect 2697 55641 2731 55675
rect 3985 55641 4019 55675
rect 5641 55641 5675 55675
rect 15209 55641 15243 55675
rect 15945 55641 15979 55675
rect 21189 55641 21223 55675
rect 25228 55641 25262 55675
rect 30205 55641 30239 55675
rect 33241 55641 33275 55675
rect 35909 55641 35943 55675
rect 37565 55641 37599 55675
rect 42625 55641 42659 55675
rect 53113 55641 53147 55675
rect 55781 55641 55815 55675
rect 56517 55641 56551 55675
rect 22109 55573 22143 55607
rect 22569 55573 22603 55607
rect 26341 55573 26375 55607
rect 28457 55573 28491 55607
rect 23213 55369 23247 55403
rect 25421 55369 25455 55403
rect 26433 55369 26467 55403
rect 36277 55369 36311 55403
rect 54677 55369 54711 55403
rect 57989 55369 58023 55403
rect 22100 55301 22134 55335
rect 57345 55301 57379 55335
rect 2329 55233 2363 55267
rect 17693 55233 17727 55267
rect 21281 55233 21315 55267
rect 21833 55233 21867 55267
rect 25605 55233 25639 55267
rect 26249 55233 26283 55267
rect 27445 55233 27479 55267
rect 27712 55233 27746 55267
rect 29469 55233 29503 55267
rect 36185 55233 36219 55267
rect 54585 55233 54619 55267
rect 55505 55233 55539 55267
rect 57897 55233 57931 55267
rect 2513 55165 2547 55199
rect 3985 55165 4019 55199
rect 17877 55165 17911 55199
rect 19257 55165 19291 55199
rect 26065 55165 26099 55199
rect 55689 55165 55723 55199
rect 29285 55097 29319 55131
rect 21097 55029 21131 55063
rect 28825 55029 28859 55063
rect 2605 54825 2639 54859
rect 3893 54825 3927 54859
rect 19349 54825 19383 54859
rect 27445 54825 27479 54859
rect 28365 54825 28399 54859
rect 28181 54689 28215 54723
rect 58173 54689 58207 54723
rect 2513 54621 2547 54655
rect 3801 54621 3835 54655
rect 19257 54621 19291 54655
rect 20085 54621 20119 54655
rect 28365 54621 28399 54655
rect 29561 54621 29595 54655
rect 56333 54621 56367 54655
rect 20352 54553 20386 54587
rect 27261 54553 27295 54587
rect 28089 54553 28123 54587
rect 29806 54553 29840 54587
rect 33241 54553 33275 54587
rect 56517 54553 56551 54587
rect 21465 54485 21499 54519
rect 27461 54485 27495 54519
rect 27629 54485 27663 54519
rect 28549 54485 28583 54519
rect 30941 54485 30975 54519
rect 33333 54485 33367 54519
rect 29653 54281 29687 54315
rect 56977 54281 57011 54315
rect 25973 54145 26007 54179
rect 26065 54145 26099 54179
rect 27905 54145 27939 54179
rect 27997 54145 28031 54179
rect 28825 54145 28859 54179
rect 28917 54145 28951 54179
rect 29837 54145 29871 54179
rect 56241 54145 56275 54179
rect 56885 54145 56919 54179
rect 58081 54145 58115 54179
rect 29009 54077 29043 54111
rect 29101 54077 29135 54111
rect 28181 54009 28215 54043
rect 26249 53941 26283 53975
rect 28641 53941 28675 53975
rect 56333 53941 56367 53975
rect 27537 53737 27571 53771
rect 28365 53737 28399 53771
rect 26985 53669 27019 53703
rect 25145 53601 25179 53635
rect 56517 53601 56551 53635
rect 58173 53601 58207 53635
rect 2237 53533 2271 53567
rect 22569 53533 22603 53567
rect 22753 53533 22787 53567
rect 27261 53533 27295 53567
rect 28595 53533 28629 53567
rect 28733 53533 28767 53567
rect 28825 53533 28859 53567
rect 29009 53533 29043 53567
rect 29561 53533 29595 53567
rect 29817 53533 29851 53567
rect 56333 53533 56367 53567
rect 25412 53465 25446 53499
rect 27353 53465 27387 53499
rect 22937 53397 22971 53431
rect 26525 53397 26559 53431
rect 27169 53397 27203 53431
rect 30941 53397 30975 53431
rect 25421 53193 25455 53227
rect 27445 53193 27479 53227
rect 1961 53057 1995 53091
rect 21833 53057 21867 53091
rect 22100 53057 22134 53091
rect 23673 53057 23707 53091
rect 23857 53057 23891 53091
rect 25605 53057 25639 53091
rect 26249 53057 26283 53091
rect 26985 53057 27019 53091
rect 27261 53057 27295 53091
rect 28089 53057 28123 53091
rect 58081 53057 58115 53091
rect 2145 52989 2179 53023
rect 2789 52989 2823 53023
rect 26065 52989 26099 53023
rect 27077 52989 27111 53023
rect 23213 52853 23247 52887
rect 24041 52853 24075 52887
rect 26433 52853 26467 52887
rect 26985 52853 27019 52887
rect 27905 52853 27939 52887
rect 2421 52649 2455 52683
rect 21465 52581 21499 52615
rect 26893 52581 26927 52615
rect 25513 52513 25547 52547
rect 2329 52445 2363 52479
rect 3157 52445 3191 52479
rect 3801 52445 3835 52479
rect 21649 52445 21683 52479
rect 22109 52445 22143 52479
rect 25780 52445 25814 52479
rect 22376 52377 22410 52411
rect 3893 52309 3927 52343
rect 23489 52309 23523 52343
rect 23305 52105 23339 52139
rect 23949 52105 23983 52139
rect 26433 52105 26467 52139
rect 26985 52105 27019 52139
rect 2421 52037 2455 52071
rect 20269 52037 20303 52071
rect 22170 52037 22204 52071
rect 24133 52037 24167 52071
rect 25320 52037 25354 52071
rect 19441 51969 19475 52003
rect 19993 51969 20027 52003
rect 20085 51969 20119 52003
rect 21925 51969 21959 52003
rect 24041 51969 24075 52003
rect 25053 51969 25087 52003
rect 27169 51969 27203 52003
rect 30205 51969 30239 52003
rect 30472 51969 30506 52003
rect 32321 51969 32355 52003
rect 32505 51969 32539 52003
rect 33149 51969 33183 52003
rect 2237 51901 2271 51935
rect 3249 51901 3283 51935
rect 32137 51901 32171 51935
rect 23765 51833 23799 51867
rect 31585 51833 31619 51867
rect 19257 51765 19291 51799
rect 24317 51765 24351 51799
rect 32965 51765 32999 51799
rect 21649 51561 21683 51595
rect 22661 51561 22695 51595
rect 23397 51561 23431 51595
rect 25973 51561 26007 51595
rect 30573 51561 30607 51595
rect 22293 51425 22327 51459
rect 23213 51425 23247 51459
rect 25605 51425 25639 51459
rect 19257 51357 19291 51391
rect 19513 51357 19547 51391
rect 21833 51357 21867 51391
rect 22477 51357 22511 51391
rect 23397 51357 23431 51391
rect 25789 51357 25823 51391
rect 29009 51357 29043 51391
rect 29745 51357 29779 51391
rect 29929 51357 29963 51391
rect 30113 51357 30147 51391
rect 30757 51357 30791 51391
rect 31309 51357 31343 51391
rect 31401 51357 31435 51391
rect 32045 51357 32079 51391
rect 32312 51357 32346 51391
rect 34069 51357 34103 51391
rect 56977 51357 57011 51391
rect 57805 51357 57839 51391
rect 23121 51289 23155 51323
rect 20637 51221 20671 51255
rect 23581 51221 23615 51255
rect 28825 51221 28859 51255
rect 31585 51221 31619 51255
rect 33425 51221 33459 51255
rect 33885 51221 33919 51255
rect 57069 51221 57103 51255
rect 23305 51017 23339 51051
rect 31585 51017 31619 51051
rect 33517 51017 33551 51051
rect 30389 50949 30423 50983
rect 30605 50949 30639 50983
rect 32404 50949 32438 50983
rect 33977 50949 34011 50983
rect 19809 50881 19843 50915
rect 19901 50881 19935 50915
rect 22569 50881 22603 50915
rect 22661 50881 22695 50915
rect 23489 50881 23523 50915
rect 24961 50881 24995 50915
rect 25697 50881 25731 50915
rect 28549 50881 28583 50915
rect 28816 50881 28850 50915
rect 31401 50881 31435 50915
rect 34253 50881 34287 50915
rect 25421 50813 25455 50847
rect 31217 50813 31251 50847
rect 32137 50813 32171 50847
rect 34069 50813 34103 50847
rect 24777 50745 24811 50779
rect 34437 50745 34471 50779
rect 20085 50677 20119 50711
rect 22845 50677 22879 50711
rect 29929 50677 29963 50711
rect 30573 50677 30607 50711
rect 30757 50677 30791 50711
rect 33977 50677 34011 50711
rect 25053 50473 25087 50507
rect 30665 50473 30699 50507
rect 33517 50473 33551 50507
rect 29009 50405 29043 50439
rect 29561 50405 29595 50439
rect 19257 50337 19291 50371
rect 26157 50337 26191 50371
rect 30849 50337 30883 50371
rect 31125 50337 31159 50371
rect 56333 50337 56367 50371
rect 56517 50337 56551 50371
rect 57897 50337 57931 50371
rect 18705 50269 18739 50303
rect 22385 50269 22419 50303
rect 25881 50269 25915 50303
rect 27629 50269 27663 50303
rect 29837 50269 29871 50303
rect 29929 50269 29963 50303
rect 30021 50269 30055 50303
rect 30205 50269 30239 50303
rect 30941 50269 30975 50303
rect 31033 50269 31067 50303
rect 32137 50269 32171 50303
rect 19502 50201 19536 50235
rect 24961 50201 24995 50235
rect 27896 50201 27930 50235
rect 32404 50201 32438 50235
rect 18521 50133 18555 50167
rect 20637 50133 20671 50167
rect 22201 50133 22235 50167
rect 18797 49929 18831 49963
rect 20453 49929 20487 49963
rect 20637 49929 20671 49963
rect 29653 49929 29687 49963
rect 30941 49929 30975 49963
rect 32321 49929 32355 49963
rect 32505 49929 32539 49963
rect 32689 49929 32723 49963
rect 33149 49929 33183 49963
rect 19809 49861 19843 49895
rect 20269 49861 20303 49895
rect 24501 49861 24535 49895
rect 27629 49861 27663 49895
rect 28540 49861 28574 49895
rect 32137 49861 32171 49895
rect 32413 49861 32447 49895
rect 18981 49793 19015 49827
rect 19625 49793 19659 49827
rect 20545 49793 20579 49827
rect 22661 49793 22695 49827
rect 23489 49793 23523 49827
rect 24317 49793 24351 49827
rect 24409 49793 24443 49827
rect 27445 49793 27479 49827
rect 28273 49793 28307 49827
rect 30297 49793 30331 49827
rect 30481 49793 30515 49827
rect 31125 49793 31159 49827
rect 33333 49793 33367 49827
rect 37832 49793 37866 49827
rect 39497 49793 39531 49827
rect 40141 49793 40175 49827
rect 40325 49793 40359 49827
rect 19441 49725 19475 49759
rect 20821 49725 20855 49759
rect 23305 49725 23339 49759
rect 23673 49725 23707 49759
rect 24685 49725 24719 49759
rect 25421 49725 25455 49759
rect 25697 49725 25731 49759
rect 30113 49725 30147 49759
rect 37565 49725 37599 49759
rect 39681 49725 39715 49759
rect 40509 49725 40543 49759
rect 24133 49657 24167 49691
rect 22477 49589 22511 49623
rect 38945 49589 38979 49623
rect 23857 49385 23891 49419
rect 29561 49385 29595 49419
rect 30021 49385 30055 49419
rect 41245 49385 41279 49419
rect 23029 49317 23063 49351
rect 29009 49317 29043 49351
rect 19257 49249 19291 49283
rect 23489 49249 23523 49283
rect 29745 49249 29779 49283
rect 39865 49249 39899 49283
rect 48973 49249 49007 49283
rect 19524 49181 19558 49215
rect 21649 49181 21683 49215
rect 21916 49181 21950 49215
rect 23673 49181 23707 49215
rect 24409 49181 24443 49215
rect 26249 49181 26283 49215
rect 26433 49181 26467 49215
rect 27629 49181 27663 49215
rect 29561 49181 29595 49215
rect 29837 49181 29871 49215
rect 30757 49181 30791 49215
rect 34713 49181 34747 49215
rect 37381 49181 37415 49215
rect 40141 49181 40175 49215
rect 41153 49181 41187 49215
rect 42073 49181 42107 49215
rect 42901 49181 42935 49215
rect 43085 49181 43119 49215
rect 47777 49181 47811 49215
rect 57069 49181 57103 49215
rect 57897 49181 57931 49215
rect 24654 49113 24688 49147
rect 27896 49113 27930 49147
rect 30573 49113 30607 49147
rect 34958 49113 34992 49147
rect 37626 49113 37660 49147
rect 42257 49113 42291 49147
rect 42441 49113 42475 49147
rect 47961 49113 47995 49147
rect 20637 49045 20671 49079
rect 25789 49045 25823 49079
rect 26617 49045 26651 49079
rect 36093 49045 36127 49079
rect 38761 49045 38795 49079
rect 41613 49045 41647 49079
rect 43177 49045 43211 49079
rect 57161 49045 57195 49079
rect 23489 48841 23523 48875
rect 26985 48841 27019 48875
rect 27813 48841 27847 48875
rect 34253 48841 34287 48875
rect 48237 48841 48271 48875
rect 20177 48773 20211 48807
rect 25320 48773 25354 48807
rect 28825 48773 28859 48807
rect 29653 48773 29687 48807
rect 33885 48773 33919 48807
rect 33977 48773 34011 48807
rect 41797 48773 41831 48807
rect 7849 48705 7883 48739
rect 20453 48705 20487 48739
rect 22109 48705 22143 48739
rect 22376 48705 22410 48739
rect 24041 48705 24075 48739
rect 24317 48705 24351 48739
rect 25053 48705 25087 48739
rect 27169 48705 27203 48739
rect 27997 48705 28031 48739
rect 28641 48705 28675 48739
rect 29469 48711 29503 48745
rect 33701 48705 33735 48739
rect 34069 48705 34103 48739
rect 37381 48705 37415 48739
rect 37648 48705 37682 48739
rect 39773 48705 39807 48739
rect 40417 48705 40451 48739
rect 41705 48705 41739 48739
rect 41889 48705 41923 48739
rect 42441 48705 42475 48739
rect 43637 48705 43671 48739
rect 43821 48705 43855 48739
rect 44741 48705 44775 48739
rect 44925 48705 44959 48739
rect 45017 48705 45051 48739
rect 45155 48705 45189 48739
rect 48145 48705 48179 48739
rect 8493 48637 8527 48671
rect 8677 48637 8711 48671
rect 9689 48637 9723 48671
rect 20269 48637 20303 48671
rect 24225 48637 24259 48671
rect 28457 48637 28491 48671
rect 29285 48637 29319 48671
rect 39221 48637 39255 48671
rect 39589 48637 39623 48671
rect 39681 48637 39715 48671
rect 40693 48637 40727 48671
rect 42625 48637 42659 48671
rect 42901 48637 42935 48671
rect 42993 48637 43027 48671
rect 7941 48569 7975 48603
rect 38761 48569 38795 48603
rect 20177 48501 20211 48535
rect 20637 48501 20671 48535
rect 24133 48501 24167 48535
rect 24501 48501 24535 48535
rect 26433 48501 26467 48535
rect 44005 48501 44039 48535
rect 45293 48501 45327 48535
rect 23673 48297 23707 48331
rect 37289 48297 37323 48331
rect 38301 48297 38335 48331
rect 46029 48297 46063 48331
rect 40141 48229 40175 48263
rect 25605 48161 25639 48195
rect 28089 48161 28123 48195
rect 41061 48161 41095 48195
rect 42533 48161 42567 48195
rect 45477 48161 45511 48195
rect 46949 48161 46983 48195
rect 56333 48161 56367 48195
rect 56517 48161 56551 48195
rect 57897 48161 57931 48195
rect 19717 48093 19751 48127
rect 19809 48093 19843 48127
rect 23857 48093 23891 48127
rect 24409 48093 24443 48127
rect 24593 48093 24627 48127
rect 25329 48093 25363 48127
rect 27813 48093 27847 48127
rect 32781 48093 32815 48127
rect 36737 48093 36771 48127
rect 37013 48093 37047 48127
rect 37105 48093 37139 48127
rect 37749 48093 37783 48127
rect 38117 48093 38151 48127
rect 39957 48093 39991 48127
rect 40601 48093 40635 48127
rect 40785 48093 40819 48127
rect 41153 48093 41187 48127
rect 42073 48093 42107 48127
rect 42257 48093 42291 48127
rect 42717 48093 42751 48127
rect 45201 48093 45235 48127
rect 45293 48093 45327 48127
rect 45569 48093 45603 48127
rect 46305 48093 46339 48127
rect 47041 48093 47075 48127
rect 47961 48093 47995 48127
rect 48145 48093 48179 48127
rect 31953 48025 31987 48059
rect 32137 48025 32171 48059
rect 33048 48025 33082 48059
rect 36921 48025 36955 48059
rect 37933 48025 37967 48059
rect 38025 48025 38059 48059
rect 44097 48025 44131 48059
rect 46029 48025 46063 48059
rect 19993 47957 20027 47991
rect 24777 47957 24811 47991
rect 32321 47957 32355 47991
rect 34161 47957 34195 47991
rect 44189 47957 44223 47991
rect 45017 47957 45051 47991
rect 46213 47957 46247 47991
rect 47409 47957 47443 47991
rect 48145 47957 48179 47991
rect 20637 47753 20671 47787
rect 33057 47753 33091 47787
rect 37841 47753 37875 47787
rect 40049 47753 40083 47787
rect 44557 47753 44591 47787
rect 46489 47753 46523 47787
rect 19064 47685 19098 47719
rect 24317 47685 24351 47719
rect 24547 47685 24581 47719
rect 25881 47685 25915 47719
rect 29745 47685 29779 47719
rect 29929 47685 29963 47719
rect 37565 47685 37599 47719
rect 40601 47685 40635 47719
rect 45017 47685 45051 47719
rect 20821 47617 20855 47651
rect 24225 47617 24259 47651
rect 24409 47617 24443 47651
rect 27445 47617 27479 47651
rect 27629 47617 27663 47651
rect 28273 47617 28307 47651
rect 30389 47617 30423 47651
rect 31125 47617 31159 47651
rect 32321 47617 32355 47651
rect 32505 47617 32539 47651
rect 32597 47617 32631 47651
rect 33333 47617 33367 47651
rect 33425 47617 33459 47651
rect 33517 47617 33551 47651
rect 33701 47617 33735 47651
rect 34161 47617 34195 47651
rect 34417 47617 34451 47651
rect 37289 47617 37323 47651
rect 37473 47617 37507 47651
rect 37657 47617 37691 47651
rect 39589 47617 39623 47651
rect 41337 47617 41371 47651
rect 41521 47617 41555 47651
rect 44189 47617 44223 47651
rect 44373 47617 44407 47651
rect 45247 47617 45281 47651
rect 45385 47617 45419 47651
rect 45477 47617 45511 47651
rect 45661 47617 45695 47651
rect 46581 47617 46615 47651
rect 47869 47617 47903 47651
rect 47958 47617 47992 47651
rect 48053 47617 48087 47651
rect 48237 47617 48271 47651
rect 48881 47617 48915 47651
rect 18797 47549 18831 47583
rect 24685 47549 24719 47583
rect 28917 47549 28951 47583
rect 46121 47549 46155 47583
rect 48789 47549 48823 47583
rect 32137 47481 32171 47515
rect 39865 47481 39899 47515
rect 46305 47481 46339 47515
rect 20177 47413 20211 47447
rect 24041 47413 24075 47447
rect 25973 47413 26007 47447
rect 30481 47413 30515 47447
rect 31217 47413 31251 47447
rect 35541 47413 35575 47447
rect 40693 47413 40727 47447
rect 41705 47413 41739 47447
rect 47593 47413 47627 47447
rect 49157 47413 49191 47447
rect 46029 47209 46063 47243
rect 47961 47209 47995 47243
rect 48237 47209 48271 47243
rect 30021 47141 30055 47175
rect 31033 47141 31067 47175
rect 19533 47073 19567 47107
rect 20729 47073 20763 47107
rect 27353 47073 27387 47107
rect 27721 47073 27755 47107
rect 30113 47073 30147 47107
rect 31677 47073 31711 47107
rect 31861 47073 31895 47107
rect 33517 47073 33551 47107
rect 46765 47073 46799 47107
rect 49157 47073 49191 47107
rect 50169 47073 50203 47107
rect 56333 47073 56367 47107
rect 19717 47005 19751 47039
rect 20361 47005 20395 47039
rect 20545 47005 20579 47039
rect 21373 47005 21407 47039
rect 22845 47005 22879 47039
rect 24409 47005 24443 47039
rect 24665 47005 24699 47039
rect 26249 47005 26283 47039
rect 27169 47005 27203 47039
rect 30849 47005 30883 47039
rect 35081 47005 35115 47039
rect 35265 47005 35299 47039
rect 36461 47005 36495 47039
rect 39957 47005 39991 47039
rect 40049 47005 40083 47039
rect 40233 47005 40267 47039
rect 40325 47005 40359 47039
rect 41429 47005 41463 47039
rect 41613 47005 41647 47039
rect 42349 47005 42383 47039
rect 44465 47005 44499 47039
rect 45201 47005 45235 47039
rect 45293 47005 45327 47039
rect 45477 47005 45511 47039
rect 45569 47005 45603 47039
rect 46305 47005 46339 47039
rect 46949 47005 46983 47039
rect 47133 47005 47167 47039
rect 47225 47005 47259 47039
rect 47685 47005 47719 47039
rect 47961 47005 47995 47039
rect 48881 47005 48915 47039
rect 48973 47005 49007 47039
rect 49249 47005 49283 47039
rect 50353 47005 50387 47039
rect 50629 47005 50663 47039
rect 19901 46937 19935 46971
rect 21189 46937 21223 46971
rect 21557 46937 21591 46971
rect 29653 46937 29687 46971
rect 35173 46937 35207 46971
rect 36277 46937 36311 46971
rect 41705 46937 41739 46971
rect 42165 46937 42199 46971
rect 42533 46937 42567 46971
rect 43085 46937 43119 46971
rect 44097 46937 44131 46971
rect 44281 46937 44315 46971
rect 46029 46937 46063 46971
rect 56517 46937 56551 46971
rect 58173 46937 58207 46971
rect 22661 46869 22695 46903
rect 25789 46869 25823 46903
rect 26433 46869 26467 46903
rect 40325 46869 40359 46903
rect 43177 46869 43211 46903
rect 45017 46869 45051 46903
rect 46213 46869 46247 46903
rect 48697 46869 48731 46903
rect 50537 46869 50571 46903
rect 24041 46665 24075 46699
rect 25605 46665 25639 46699
rect 27629 46665 27663 46699
rect 31401 46665 31435 46699
rect 42625 46665 42659 46699
rect 45109 46665 45143 46699
rect 51089 46665 51123 46699
rect 56977 46665 57011 46699
rect 19340 46597 19374 46631
rect 22201 46597 22235 46631
rect 22319 46597 22353 46631
rect 23029 46597 23063 46631
rect 26249 46597 26283 46631
rect 27537 46597 27571 46631
rect 44741 46597 44775 46631
rect 44957 46597 44991 46631
rect 19073 46529 19107 46563
rect 22017 46529 22051 46563
rect 22109 46529 22143 46563
rect 22477 46529 22511 46563
rect 23857 46529 23891 46563
rect 24777 46529 24811 46563
rect 25513 46529 25547 46563
rect 28273 46529 28307 46563
rect 30021 46529 30055 46563
rect 30288 46529 30322 46563
rect 32413 46529 32447 46563
rect 32502 46529 32536 46563
rect 32597 46532 32631 46566
rect 32781 46529 32815 46563
rect 34161 46529 34195 46563
rect 36093 46529 36127 46563
rect 37933 46529 37967 46563
rect 38117 46529 38151 46563
rect 39221 46529 39255 46563
rect 39405 46529 39439 46563
rect 40141 46529 40175 46563
rect 40230 46535 40264 46569
rect 40325 46529 40359 46563
rect 40509 46529 40543 46563
rect 42441 46529 42475 46563
rect 42717 46529 42751 46563
rect 43361 46529 43395 46563
rect 43545 46529 43579 46563
rect 43637 46529 43671 46563
rect 43913 46529 43947 46563
rect 45569 46529 45603 46563
rect 45753 46529 45787 46563
rect 46857 46529 46891 46563
rect 49893 46529 49927 46563
rect 50077 46529 50111 46563
rect 50721 46529 50755 46563
rect 56885 46529 56919 46563
rect 58081 46529 58115 46563
rect 23673 46461 23707 46495
rect 24593 46461 24627 46495
rect 29377 46461 29411 46495
rect 34437 46461 34471 46495
rect 35817 46461 35851 46495
rect 43729 46461 43763 46495
rect 45661 46461 45695 46495
rect 47593 46461 47627 46495
rect 47869 46461 47903 46495
rect 50813 46461 50847 46495
rect 26433 46393 26467 46427
rect 39865 46393 39899 46427
rect 20453 46325 20487 46359
rect 21833 46325 21867 46359
rect 23121 46325 23155 46359
rect 24961 46325 24995 46359
rect 32137 46325 32171 46359
rect 38025 46325 38059 46359
rect 39221 46325 39255 46359
rect 42441 46325 42475 46359
rect 44097 46325 44131 46359
rect 44925 46325 44959 46359
rect 46949 46325 46983 46359
rect 49893 46325 49927 46359
rect 20637 46121 20671 46155
rect 27077 46121 27111 46155
rect 29009 46121 29043 46155
rect 34805 46121 34839 46155
rect 45109 46121 45143 46155
rect 45661 46121 45695 46155
rect 47777 46121 47811 46155
rect 47961 46121 47995 46155
rect 21097 46053 21131 46087
rect 23121 46053 23155 46087
rect 18337 45985 18371 46019
rect 19257 45985 19291 46019
rect 21741 45985 21775 46019
rect 24409 45985 24443 46019
rect 29929 45985 29963 46019
rect 31033 45985 31067 46019
rect 36277 45985 36311 46019
rect 18521 45917 18555 45951
rect 21281 45917 21315 45951
rect 23857 45917 23891 45951
rect 27629 45917 27663 45951
rect 29561 45917 29595 45951
rect 31300 45917 31334 45951
rect 33425 45917 33459 45951
rect 33517 45917 33551 45951
rect 33609 45917 33643 45951
rect 33793 45917 33827 45951
rect 34713 45917 34747 45951
rect 34897 45917 34931 45951
rect 36001 45917 36035 45951
rect 36093 45917 36127 45951
rect 37657 45917 37691 45951
rect 37933 45917 37967 45951
rect 38117 45917 38151 45951
rect 38577 45917 38611 45951
rect 38945 45917 38979 45951
rect 40141 45917 40175 45951
rect 40233 45917 40267 45951
rect 40325 45917 40359 45951
rect 40509 45917 40543 45951
rect 41061 45917 41095 45951
rect 41245 45917 41279 45951
rect 42349 45917 42383 45951
rect 42717 45917 42751 45951
rect 42809 45917 42843 45951
rect 44189 45917 44223 45951
rect 45017 45917 45051 45951
rect 45201 45917 45235 45951
rect 45661 45917 45695 45951
rect 45845 45917 45879 45951
rect 50997 45917 51031 45951
rect 51273 45917 51307 45951
rect 56977 45917 57011 45951
rect 57805 45917 57839 45951
rect 19502 45849 19536 45883
rect 21986 45849 22020 45883
rect 24676 45849 24710 45883
rect 26985 45849 27019 45883
rect 27874 45849 27908 45883
rect 38761 45849 38795 45883
rect 38853 45849 38887 45883
rect 42441 45849 42475 45883
rect 42533 45849 42567 45883
rect 47593 45849 47627 45883
rect 50813 45849 50847 45883
rect 18705 45781 18739 45815
rect 23673 45781 23707 45815
rect 25789 45781 25823 45815
rect 32413 45781 32447 45815
rect 33149 45781 33183 45815
rect 36277 45781 36311 45815
rect 37841 45781 37875 45815
rect 39129 45781 39163 45815
rect 39865 45781 39899 45815
rect 41153 45781 41187 45815
rect 42165 45781 42199 45815
rect 44281 45781 44315 45815
rect 47793 45781 47827 45815
rect 51181 45781 51215 45815
rect 57069 45781 57103 45815
rect 21005 45577 21039 45611
rect 34437 45577 34471 45611
rect 38945 45577 38979 45611
rect 48053 45577 48087 45611
rect 22652 45509 22686 45543
rect 25145 45509 25179 45543
rect 27353 45509 27387 45543
rect 27997 45509 28031 45543
rect 30113 45509 30147 45543
rect 32404 45509 32438 45543
rect 40233 45509 40267 45543
rect 45753 45509 45787 45543
rect 49433 45509 49467 45543
rect 53205 45509 53239 45543
rect 55781 45509 55815 45543
rect 18889 45441 18923 45475
rect 19156 45441 19190 45475
rect 20729 45441 20763 45475
rect 20913 45441 20947 45475
rect 21097 45441 21131 45475
rect 21281 45441 21315 45475
rect 26065 45441 26099 45475
rect 26249 45441 26283 45475
rect 27721 45441 27755 45475
rect 28273 45441 28307 45475
rect 34345 45441 34379 45475
rect 34529 45441 34563 45475
rect 34989 45441 35023 45475
rect 35173 45441 35207 45475
rect 35357 45441 35391 45475
rect 35541 45441 35575 45475
rect 36461 45441 36495 45475
rect 36645 45441 36679 45475
rect 36737 45441 36771 45475
rect 37565 45441 37599 45475
rect 37749 45441 37783 45475
rect 37842 45441 37876 45475
rect 38577 45441 38611 45475
rect 40417 45441 40451 45475
rect 40509 45441 40543 45475
rect 40693 45441 40727 45475
rect 40877 45441 40911 45475
rect 41705 45441 41739 45475
rect 41797 45441 41831 45475
rect 42441 45441 42475 45475
rect 42625 45441 42659 45475
rect 42717 45441 42751 45475
rect 42993 45441 43027 45475
rect 45937 45441 45971 45475
rect 46029 45441 46063 45475
rect 46765 45441 46799 45475
rect 47593 45441 47627 45475
rect 47869 45441 47903 45475
rect 48605 45441 48639 45475
rect 48973 45441 49007 45475
rect 49157 45441 49191 45475
rect 51457 45441 51491 45475
rect 55965 45441 55999 45475
rect 56057 45441 56091 45475
rect 22385 45373 22419 45407
rect 24225 45373 24259 45407
rect 29009 45373 29043 45407
rect 32137 45373 32171 45407
rect 35265 45373 35299 45407
rect 37646 45373 37680 45407
rect 38669 45373 38703 45407
rect 41521 45373 41555 45407
rect 41613 45373 41647 45407
rect 42809 45373 42843 45407
rect 47685 45373 47719 45407
rect 51549 45373 51583 45407
rect 51825 45373 51859 45407
rect 23765 45305 23799 45339
rect 24593 45305 24627 45339
rect 25421 45305 25455 45339
rect 30297 45305 30331 45339
rect 40601 45305 40635 45339
rect 43177 45305 43211 45339
rect 49065 45305 49099 45339
rect 20269 45237 20303 45271
rect 24685 45237 24719 45271
rect 25605 45237 25639 45271
rect 26065 45237 26099 45271
rect 33517 45237 33551 45271
rect 35725 45237 35759 45271
rect 36461 45237 36495 45271
rect 37381 45237 37415 45271
rect 41337 45237 41371 45271
rect 45753 45237 45787 45271
rect 46857 45237 46891 45271
rect 47593 45237 47627 45271
rect 53297 45237 53331 45271
rect 55781 45237 55815 45271
rect 19257 45033 19291 45067
rect 20177 45033 20211 45067
rect 20545 45033 20579 45067
rect 24961 45033 24995 45067
rect 27353 45033 27387 45067
rect 38393 45033 38427 45067
rect 39129 45033 39163 45067
rect 40325 45033 40359 45067
rect 46581 45033 46615 45067
rect 46949 45033 46983 45067
rect 48145 45033 48179 45067
rect 49617 45033 49651 45067
rect 53481 45033 53515 45067
rect 37105 44965 37139 44999
rect 38669 44965 38703 44999
rect 55505 44965 55539 44999
rect 20269 44897 20303 44931
rect 25881 44897 25915 44931
rect 29929 44897 29963 44931
rect 30757 44897 30791 44931
rect 37289 44897 37323 44931
rect 37381 44897 37415 44931
rect 49249 44897 49283 44931
rect 56333 44897 56367 44931
rect 56517 44897 56551 44931
rect 57897 44897 57931 44931
rect 19441 44829 19475 44863
rect 20361 44829 20395 44863
rect 24685 44829 24719 44863
rect 24777 44829 24811 44863
rect 25053 44829 25087 44863
rect 25605 44829 25639 44863
rect 25697 44829 25731 44863
rect 27537 44829 27571 44863
rect 28181 44829 28215 44863
rect 29561 44829 29595 44863
rect 29745 44829 29779 44863
rect 32827 44829 32861 44863
rect 32965 44829 32999 44863
rect 33057 44829 33091 44863
rect 33241 44829 33275 44863
rect 34713 44829 34747 44863
rect 34980 44829 35014 44863
rect 37473 44829 37507 44863
rect 37565 44829 37599 44863
rect 38117 44829 38151 44863
rect 38393 44829 38427 44863
rect 39129 44829 39163 44863
rect 39313 44829 39347 44863
rect 40509 44829 40543 44863
rect 40877 44829 40911 44863
rect 40969 44829 41003 44863
rect 42165 44829 42199 44863
rect 42441 44829 42475 44863
rect 43269 44829 43303 44863
rect 45477 44829 45511 44863
rect 46489 44829 46523 44863
rect 47777 44829 47811 44863
rect 47961 44829 47995 44863
rect 49433 44829 49467 44863
rect 50721 44829 50755 44863
rect 50997 44829 51031 44863
rect 51457 44829 51491 44863
rect 51641 44829 51675 44863
rect 51917 44829 51951 44863
rect 52101 44829 52135 44863
rect 52745 44829 52779 44863
rect 53021 44829 53055 44863
rect 53481 44829 53515 44863
rect 53665 44829 53699 44863
rect 55505 44829 55539 44863
rect 55689 44829 55723 44863
rect 55873 44829 55907 44863
rect 20085 44761 20119 44795
rect 28825 44761 28859 44795
rect 31024 44761 31058 44795
rect 32597 44761 32631 44795
rect 40601 44761 40635 44795
rect 40693 44761 40727 44795
rect 42901 44761 42935 44795
rect 43085 44761 43119 44795
rect 52561 44761 52595 44795
rect 24501 44693 24535 44727
rect 32137 44693 32171 44727
rect 36093 44693 36127 44727
rect 41981 44693 42015 44727
rect 42349 44693 42383 44727
rect 45569 44693 45603 44727
rect 50537 44693 50571 44727
rect 50905 44693 50939 44727
rect 52929 44693 52963 44727
rect 19533 44489 19567 44523
rect 39697 44489 39731 44523
rect 39865 44489 39899 44523
rect 43729 44489 43763 44523
rect 48237 44489 48271 44523
rect 49249 44489 49283 44523
rect 52101 44489 52135 44523
rect 53665 44489 53699 44523
rect 33784 44421 33818 44455
rect 35357 44421 35391 44455
rect 39497 44421 39531 44455
rect 41429 44421 41463 44455
rect 45569 44421 45603 44455
rect 50169 44421 50203 44455
rect 50997 44421 51031 44455
rect 51181 44421 51215 44455
rect 54493 44421 54527 44455
rect 54677 44421 54711 44455
rect 55229 44421 55263 44455
rect 55873 44421 55907 44455
rect 56701 44421 56735 44455
rect 19717 44353 19751 44387
rect 24685 44353 24719 44387
rect 24777 44353 24811 44387
rect 25053 44353 25087 44387
rect 28089 44353 28123 44387
rect 28356 44353 28390 44387
rect 32413 44353 32447 44387
rect 32505 44353 32539 44387
rect 32597 44353 32631 44387
rect 32781 44353 32815 44387
rect 33517 44353 33551 44387
rect 35633 44353 35667 44387
rect 35725 44353 35759 44387
rect 35817 44353 35851 44387
rect 36001 44353 36035 44387
rect 41337 44353 41371 44387
rect 42625 44353 42659 44387
rect 42717 44353 42751 44387
rect 42901 44353 42935 44387
rect 42993 44353 43027 44387
rect 43453 44353 43487 44387
rect 44833 44353 44867 44387
rect 45017 44353 45051 44387
rect 46490 44353 46524 44387
rect 46673 44353 46707 44387
rect 47869 44353 47903 44387
rect 48053 44353 48087 44387
rect 49157 44353 49191 44387
rect 49341 44353 49375 44387
rect 50077 44353 50111 44387
rect 50261 44353 50295 44387
rect 50813 44353 50847 44387
rect 52009 44353 52043 44387
rect 52193 44353 52227 44387
rect 52745 44353 52779 44387
rect 52929 44353 52963 44387
rect 53573 44353 53607 44387
rect 53757 44353 53791 44387
rect 54769 44353 54803 44387
rect 55689 44353 55723 44387
rect 56517 44353 56551 44387
rect 56793 44353 56827 44387
rect 43545 44285 43579 44319
rect 43729 44285 43763 44319
rect 46397 44285 46431 44319
rect 46582 44285 46616 44319
rect 55597 44285 55631 44319
rect 56333 44285 56367 44319
rect 24961 44217 24995 44251
rect 45753 44217 45787 44251
rect 24501 44149 24535 44183
rect 29469 44149 29503 44183
rect 32137 44149 32171 44183
rect 34897 44149 34931 44183
rect 39681 44149 39715 44183
rect 42441 44149 42475 44183
rect 44925 44149 44959 44183
rect 46213 44149 46247 44183
rect 53113 44149 53147 44183
rect 54493 44149 54527 44183
rect 58081 44149 58115 44183
rect 29561 43945 29595 43979
rect 35771 43945 35805 43979
rect 37749 43945 37783 43979
rect 39865 43945 39899 43979
rect 43085 43945 43119 43979
rect 50169 43945 50203 43979
rect 52653 43945 52687 43979
rect 53849 43945 53883 43979
rect 55505 43945 55539 43979
rect 39221 43877 39255 43911
rect 42533 43877 42567 43911
rect 47501 43877 47535 43911
rect 47593 43877 47627 43911
rect 48237 43877 48271 43911
rect 55689 43877 55723 43911
rect 27813 43809 27847 43843
rect 31125 43809 31159 43843
rect 38209 43809 38243 43843
rect 38853 43809 38887 43843
rect 40325 43809 40359 43843
rect 45201 43809 45235 43843
rect 46673 43809 46707 43843
rect 46765 43809 46799 43843
rect 50721 43809 50755 43843
rect 52377 43809 52411 43843
rect 56333 43809 56367 43843
rect 57897 43809 57931 43843
rect 27997 43741 28031 43775
rect 28181 43741 28215 43775
rect 29745 43741 29779 43775
rect 31392 43741 31426 43775
rect 35541 43741 35575 43775
rect 37933 43741 37967 43775
rect 38025 43741 38059 43775
rect 38117 43741 38151 43775
rect 38761 43741 38795 43775
rect 38945 43741 38979 43775
rect 39037 43741 39071 43775
rect 39313 43741 39347 43775
rect 40049 43741 40083 43775
rect 40141 43741 40175 43775
rect 40417 43741 40451 43775
rect 41337 43741 41371 43775
rect 41429 43741 41463 43775
rect 41613 43741 41647 43775
rect 41715 43741 41749 43775
rect 44097 43741 44131 43775
rect 44189 43741 44223 43775
rect 44373 43741 44407 43775
rect 44465 43741 44499 43775
rect 45293 43741 45327 43775
rect 46305 43741 46339 43775
rect 46397 43741 46431 43775
rect 47409 43741 47443 43775
rect 47685 43741 47719 43775
rect 48237 43741 48271 43775
rect 48421 43741 48455 43775
rect 50350 43741 50384 43775
rect 50813 43741 50847 43775
rect 52285 43741 52319 43775
rect 53757 43741 53791 43775
rect 53941 43741 53975 43775
rect 54401 43741 54435 43775
rect 54585 43741 54619 43775
rect 42809 43673 42843 43707
rect 43913 43673 43947 43707
rect 45569 43673 45603 43707
rect 45661 43673 45695 43707
rect 55321 43673 55355 43707
rect 56517 43673 56551 43707
rect 32505 43605 32539 43639
rect 41153 43605 41187 43639
rect 42717 43605 42751 43639
rect 42901 43605 42935 43639
rect 45017 43605 45051 43639
rect 46121 43605 46155 43639
rect 47225 43605 47259 43639
rect 50353 43605 50387 43639
rect 54769 43605 54803 43639
rect 55521 43605 55555 43639
rect 25513 43401 25547 43435
rect 41337 43401 41371 43435
rect 43177 43401 43211 43435
rect 43729 43401 43763 43435
rect 44741 43401 44775 43435
rect 46029 43401 46063 43435
rect 46489 43401 46523 43435
rect 50721 43401 50755 43435
rect 51641 43401 51675 43435
rect 54309 43401 54343 43435
rect 55137 43401 55171 43435
rect 55505 43401 55539 43435
rect 57161 43401 57195 43435
rect 25329 43333 25363 43367
rect 38669 43333 38703 43367
rect 43821 43333 43855 43367
rect 44373 43333 44407 43367
rect 47869 43333 47903 43367
rect 22293 43265 22327 43299
rect 23121 43265 23155 43299
rect 24133 43265 24167 43299
rect 26157 43265 26191 43299
rect 26341 43265 26375 43299
rect 26433 43265 26467 43299
rect 34805 43265 34839 43299
rect 34989 43265 35023 43299
rect 35081 43265 35115 43299
rect 35357 43265 35391 43299
rect 36001 43265 36035 43299
rect 36185 43265 36219 43299
rect 36277 43265 36311 43299
rect 36553 43265 36587 43299
rect 38393 43265 38427 43299
rect 41245 43265 41279 43299
rect 41429 43265 41463 43299
rect 42441 43265 42475 43299
rect 42625 43265 42659 43299
rect 42717 43265 42751 43299
rect 42993 43265 43027 43299
rect 43637 43265 43671 43299
rect 43913 43265 43947 43299
rect 44557 43265 44591 43299
rect 44833 43265 44867 43299
rect 45293 43265 45327 43299
rect 45477 43265 45511 43299
rect 45569 43265 45603 43299
rect 45845 43265 45879 43299
rect 46673 43265 46707 43299
rect 47593 43265 47627 43299
rect 47685 43265 47719 43299
rect 49065 43265 49099 43299
rect 50838 43265 50872 43299
rect 51457 43265 51491 43299
rect 52745 43265 52779 43299
rect 52929 43265 52963 43299
rect 53205 43265 53239 43299
rect 53481 43265 53515 43299
rect 54217 43265 54251 43299
rect 54401 43265 54435 43299
rect 55321 43265 55355 43299
rect 55597 43265 55631 43299
rect 56333 43265 56367 43299
rect 57897 43265 57931 43299
rect 24225 43197 24259 43231
rect 24317 43197 24351 43231
rect 24409 43197 24443 43231
rect 35173 43197 35207 43231
rect 36369 43197 36403 43231
rect 38669 43197 38703 43231
rect 40969 43197 41003 43231
rect 41705 43197 41739 43231
rect 42809 43197 42843 43231
rect 45661 43197 45695 43231
rect 46857 43197 46891 43231
rect 46949 43197 46983 43231
rect 47869 43197 47903 43231
rect 49341 43197 49375 43231
rect 50353 43197 50387 43231
rect 50629 43197 50663 43231
rect 56517 43197 56551 43231
rect 24961 43129 24995 43163
rect 50997 43129 51031 43163
rect 53113 43129 53147 43163
rect 22569 43061 22603 43095
rect 23305 43061 23339 43095
rect 23949 43061 23983 43095
rect 25329 43061 25363 43095
rect 25973 43061 26007 43095
rect 35541 43061 35575 43095
rect 36737 43061 36771 43095
rect 38485 43061 38519 43095
rect 41613 43061 41647 43095
rect 57989 43061 58023 43095
rect 37749 42857 37783 42891
rect 38761 42857 38795 42891
rect 41337 42857 41371 42891
rect 42625 42857 42659 42891
rect 46673 42857 46707 42891
rect 48237 42857 48271 42891
rect 51365 42857 51399 42891
rect 53113 42857 53147 42891
rect 55413 42857 55447 42891
rect 22569 42789 22603 42823
rect 23581 42789 23615 42823
rect 23673 42789 23707 42823
rect 41889 42789 41923 42823
rect 20361 42721 20395 42755
rect 20637 42721 20671 42755
rect 25329 42721 25363 42755
rect 30573 42721 30607 42755
rect 31953 42721 31987 42755
rect 32689 42721 32723 42755
rect 37565 42721 37599 42755
rect 38393 42721 38427 42755
rect 41981 42721 42015 42755
rect 45753 42721 45787 42755
rect 47225 42721 47259 42755
rect 52837 42721 52871 42755
rect 54401 42721 54435 42755
rect 56517 42721 56551 42755
rect 57897 42721 57931 42755
rect 20269 42653 20303 42687
rect 21189 42653 21223 42687
rect 23489 42653 23523 42687
rect 23765 42653 23799 42687
rect 24409 42653 24443 42687
rect 24685 42653 24719 42687
rect 28273 42653 28307 42687
rect 29745 42653 29779 42687
rect 30205 42653 30239 42687
rect 30389 42653 30423 42687
rect 31585 42653 31619 42687
rect 31769 42653 31803 42687
rect 32505 42653 32539 42687
rect 34713 42653 34747 42687
rect 34980 42653 35014 42687
rect 37473 42653 37507 42687
rect 38485 42653 38519 42687
rect 41462 42653 41496 42687
rect 42441 42653 42475 42687
rect 42625 42653 42659 42687
rect 45017 42653 45051 42687
rect 45201 42653 45235 42687
rect 45293 42653 45327 42687
rect 45385 42653 45419 42687
rect 45569 42653 45603 42687
rect 46305 42653 46339 42687
rect 47133 42653 47167 42687
rect 47317 42653 47351 42687
rect 48145 42653 48179 42687
rect 48329 42653 48363 42687
rect 51273 42653 51307 42687
rect 51457 42653 51491 42687
rect 52745 42653 52779 42687
rect 55597 42653 55631 42687
rect 56333 42653 56367 42687
rect 21434 42585 21468 42619
rect 23305 42585 23339 42619
rect 25596 42585 25630 42619
rect 27261 42585 27295 42619
rect 27445 42585 27479 42619
rect 46489 42585 46523 42619
rect 50629 42585 50663 42619
rect 54033 42585 54067 42619
rect 54217 42585 54251 42619
rect 55321 42585 55355 42619
rect 55505 42585 55539 42619
rect 24507 42517 24541 42551
rect 24593 42517 24627 42551
rect 26709 42517 26743 42551
rect 28089 42517 28123 42551
rect 29561 42517 29595 42551
rect 36093 42517 36127 42551
rect 41521 42517 41555 42551
rect 42809 42517 42843 42551
rect 50721 42517 50755 42551
rect 20913 42313 20947 42347
rect 25237 42313 25271 42347
rect 25789 42313 25823 42347
rect 29561 42313 29595 42347
rect 35633 42313 35667 42347
rect 38669 42313 38703 42347
rect 41711 42313 41745 42347
rect 42809 42313 42843 42347
rect 50077 42313 50111 42347
rect 51825 42313 51859 42347
rect 54493 42313 54527 42347
rect 55413 42313 55447 42347
rect 56977 42313 57011 42347
rect 32413 42245 32447 42279
rect 39313 42245 39347 42279
rect 41613 42245 41647 42279
rect 42441 42245 42475 42279
rect 48605 42245 48639 42279
rect 42671 42211 42705 42245
rect 19533 42177 19567 42211
rect 19800 42177 19834 42211
rect 22017 42177 22051 42211
rect 23857 42177 23891 42211
rect 24113 42177 24147 42211
rect 25973 42177 26007 42211
rect 26249 42177 26283 42211
rect 26433 42177 26467 42211
rect 27537 42177 27571 42211
rect 28273 42177 28307 42211
rect 30665 42177 30699 42211
rect 31217 42177 31251 42211
rect 31401 42177 31435 42211
rect 32137 42177 32171 42211
rect 32321 42177 32355 42211
rect 32505 42177 32539 42211
rect 34253 42177 34287 42211
rect 34520 42177 34554 42211
rect 38301 42177 38335 42211
rect 39129 42177 39163 42211
rect 40509 42177 40543 42211
rect 40693 42177 40727 42211
rect 41797 42177 41831 42211
rect 41889 42177 41923 42211
rect 43269 42177 43303 42211
rect 43453 42177 43487 42211
rect 47777 42177 47811 42211
rect 47869 42177 47903 42211
rect 48513 42177 48547 42211
rect 48697 42177 48731 42211
rect 49985 42177 50019 42211
rect 50169 42177 50203 42211
rect 51733 42177 51767 42211
rect 51917 42177 51951 42211
rect 54125 42177 54159 42211
rect 54953 42177 54987 42211
rect 56885 42177 56919 42211
rect 57069 42177 57103 42211
rect 58081 42177 58115 42211
rect 21925 42109 21959 42143
rect 38393 42109 38427 42143
rect 39497 42109 39531 42143
rect 54217 42109 54251 42143
rect 32689 42041 32723 42075
rect 43269 42041 43303 42075
rect 48053 42041 48087 42075
rect 22293 41973 22327 42007
rect 27721 41973 27755 42007
rect 30481 41973 30515 42007
rect 31217 41973 31251 42007
rect 40785 41973 40819 42007
rect 42625 41973 42659 42007
rect 55045 41973 55079 42007
rect 20177 41769 20211 41803
rect 21281 41769 21315 41803
rect 22385 41769 22419 41803
rect 23581 41769 23615 41803
rect 24961 41769 24995 41803
rect 28089 41769 28123 41803
rect 29009 41769 29043 41803
rect 31493 41769 31527 41803
rect 33057 41769 33091 41803
rect 37105 41769 37139 41803
rect 42441 41769 42475 41803
rect 48605 41769 48639 41803
rect 56701 41769 56735 41803
rect 28917 41701 28951 41735
rect 47869 41701 47903 41735
rect 27721 41633 27755 41667
rect 28549 41633 28583 41667
rect 32597 41633 32631 41667
rect 38025 41633 38059 41667
rect 19533 41565 19567 41599
rect 19717 41565 19751 41599
rect 20453 41565 20487 41599
rect 20545 41565 20579 41599
rect 20658 41565 20692 41599
rect 20821 41565 20855 41599
rect 21511 41565 21545 41599
rect 21646 41565 21680 41599
rect 21746 41565 21780 41599
rect 21925 41565 21959 41599
rect 22569 41565 22603 41599
rect 22845 41565 22879 41599
rect 23857 41565 23891 41599
rect 24869 41565 24903 41599
rect 27077 41565 27111 41599
rect 27905 41565 27939 41599
rect 30113 41565 30147 41599
rect 30369 41565 30403 41599
rect 32137 41565 32171 41599
rect 32322 41565 32356 41599
rect 33241 41565 33275 41599
rect 33517 41565 33551 41599
rect 37289 41565 37323 41599
rect 37565 41565 37599 41599
rect 38209 41565 38243 41599
rect 38485 41565 38519 41599
rect 38669 41565 38703 41599
rect 42441 41565 42475 41599
rect 42625 41565 42659 41599
rect 45109 41565 45143 41599
rect 45201 41565 45235 41599
rect 48421 41565 48455 41599
rect 50721 41565 50755 41599
rect 51181 41565 51215 41599
rect 51365 41565 51399 41599
rect 56977 41565 57011 41599
rect 22753 41497 22787 41531
rect 23581 41497 23615 41531
rect 32229 41497 32263 41531
rect 32439 41497 32473 41531
rect 47501 41497 47535 41531
rect 56701 41497 56735 41531
rect 19625 41429 19659 41463
rect 23765 41429 23799 41463
rect 27169 41429 27203 41463
rect 31953 41429 31987 41463
rect 33425 41429 33459 41463
rect 37473 41429 37507 41463
rect 45293 41429 45327 41463
rect 47961 41429 47995 41463
rect 50537 41429 50571 41463
rect 51365 41429 51399 41463
rect 56885 41429 56919 41463
rect 22201 41225 22235 41259
rect 24133 41225 24167 41259
rect 33517 41225 33551 41259
rect 34069 41225 34103 41259
rect 38301 41225 38335 41259
rect 39221 41225 39255 41259
rect 40049 41225 40083 41259
rect 41613 41225 41647 41259
rect 43177 41225 43211 41259
rect 49249 41225 49283 41259
rect 49893 41225 49927 41259
rect 50077 41225 50111 41259
rect 51273 41225 51307 41259
rect 51549 41225 51583 41259
rect 56333 41225 56367 41259
rect 57253 41225 57287 41259
rect 32321 41157 32355 41191
rect 32413 41157 32447 41191
rect 39681 41157 39715 41191
rect 48053 41157 48087 41191
rect 48881 41157 48915 41191
rect 56885 41157 56919 41191
rect 57101 41157 57135 41191
rect 20637 41089 20671 41123
rect 22017 41089 22051 41123
rect 23949 41089 23983 41123
rect 24133 41089 24167 41123
rect 24593 41089 24627 41123
rect 27905 41089 27939 41123
rect 29653 41089 29687 41123
rect 29837 41089 29871 41123
rect 30297 41089 30331 41123
rect 30573 41089 30607 41123
rect 32137 41089 32171 41123
rect 32505 41089 32539 41123
rect 33149 41089 33183 41123
rect 33333 41089 33367 41123
rect 33977 41089 34011 41123
rect 34161 41089 34195 41123
rect 38025 41089 38059 41123
rect 38301 41089 38335 41123
rect 39037 41089 39071 41123
rect 39865 41089 39899 41123
rect 40601 41089 40635 41123
rect 40785 41089 40819 41123
rect 41521 41089 41555 41123
rect 41705 41089 41739 41123
rect 42901 41089 42935 41123
rect 42993 41089 43027 41123
rect 46857 41089 46891 41123
rect 47777 41089 47811 41123
rect 47870 41089 47904 41123
rect 48145 41089 48179 41123
rect 48242 41089 48276 41123
rect 49065 41089 49099 41123
rect 50074 41089 50108 41123
rect 50997 41089 51031 41123
rect 51181 41089 51215 41123
rect 51365 41089 51399 41123
rect 52009 41089 52043 41123
rect 52193 41089 52227 41123
rect 56241 41089 56275 41123
rect 56425 41089 56459 41123
rect 20545 41021 20579 41055
rect 21005 41021 21039 41055
rect 21833 41021 21867 41055
rect 24869 41021 24903 41055
rect 27629 41021 27663 41055
rect 38853 41021 38887 41055
rect 50537 41021 50571 41055
rect 24777 40953 24811 40987
rect 24685 40885 24719 40919
rect 28641 40885 28675 40919
rect 29653 40885 29687 40919
rect 32689 40885 32723 40919
rect 40601 40885 40635 40919
rect 46949 40885 46983 40919
rect 48421 40885 48455 40919
rect 50445 40885 50479 40919
rect 52101 40885 52135 40919
rect 57069 40885 57103 40919
rect 21097 40681 21131 40715
rect 21189 40681 21223 40715
rect 21833 40681 21867 40715
rect 29929 40681 29963 40715
rect 31309 40681 31343 40715
rect 31493 40681 31527 40715
rect 35081 40681 35115 40715
rect 37013 40681 37047 40715
rect 42165 40681 42199 40715
rect 47225 40681 47259 40715
rect 48421 40681 48455 40715
rect 49525 40681 49559 40715
rect 56701 40681 56735 40715
rect 57253 40681 57287 40715
rect 24409 40613 24443 40647
rect 33517 40613 33551 40647
rect 39865 40613 39899 40647
rect 50445 40613 50479 40647
rect 21281 40545 21315 40579
rect 24777 40545 24811 40579
rect 28181 40545 28215 40579
rect 30481 40545 30515 40579
rect 31953 40545 31987 40579
rect 38853 40545 38887 40579
rect 40049 40545 40083 40579
rect 40417 40545 40451 40579
rect 43085 40545 43119 40579
rect 46581 40545 46615 40579
rect 51641 40545 51675 40579
rect 21005 40477 21039 40511
rect 21741 40477 21775 40511
rect 21925 40477 21959 40511
rect 24593 40477 24627 40511
rect 24869 40477 24903 40511
rect 27721 40477 27755 40511
rect 28365 40477 28399 40511
rect 30389 40477 30423 40511
rect 32229 40477 32263 40511
rect 33333 40477 33367 40511
rect 34897 40477 34931 40511
rect 35173 40477 35207 40511
rect 37013 40477 37047 40511
rect 37197 40477 37231 40511
rect 38577 40477 38611 40511
rect 38761 40477 38795 40511
rect 38945 40477 38979 40511
rect 39129 40477 39163 40511
rect 40141 40477 40175 40511
rect 41061 40477 41095 40511
rect 41245 40477 41279 40511
rect 41521 40477 41555 40511
rect 41717 40477 41751 40511
rect 42165 40477 42199 40511
rect 42349 40477 42383 40511
rect 42901 40477 42935 40511
rect 46709 40471 46743 40505
rect 47409 40477 47443 40511
rect 47593 40477 47627 40511
rect 47869 40477 47903 40511
rect 48329 40477 48363 40511
rect 48513 40477 48547 40511
rect 50169 40477 50203 40511
rect 50353 40477 50387 40511
rect 51549 40477 51583 40511
rect 52377 40477 52411 40511
rect 55505 40477 55539 40511
rect 55781 40477 55815 40511
rect 56333 40477 56367 40511
rect 57161 40477 57195 40511
rect 57345 40477 57379 40511
rect 23213 40409 23247 40443
rect 25329 40409 25363 40443
rect 25513 40409 25547 40443
rect 28549 40409 28583 40443
rect 31125 40409 31159 40443
rect 40509 40409 40543 40443
rect 46305 40409 46339 40443
rect 46489 40409 46523 40443
rect 46581 40409 46615 40443
rect 47501 40409 47535 40443
rect 47711 40409 47745 40443
rect 49433 40409 49467 40443
rect 55689 40409 55723 40443
rect 56517 40409 56551 40443
rect 23305 40341 23339 40375
rect 25697 40341 25731 40375
rect 27537 40341 27571 40375
rect 30297 40341 30331 40375
rect 31325 40341 31359 40375
rect 34713 40341 34747 40375
rect 39313 40341 39347 40375
rect 51917 40341 51951 40375
rect 52561 40341 52595 40375
rect 55321 40341 55355 40375
rect 23949 40137 23983 40171
rect 25789 40137 25823 40171
rect 30113 40137 30147 40171
rect 37933 40137 37967 40171
rect 38485 40137 38519 40171
rect 40969 40137 41003 40171
rect 51457 40137 51491 40171
rect 51641 40137 51675 40171
rect 56517 40137 56551 40171
rect 22293 40069 22327 40103
rect 30021 40069 30055 40103
rect 32229 40069 32263 40103
rect 33149 40069 33183 40103
rect 33249 40069 33283 40103
rect 39497 40069 39531 40103
rect 40601 40069 40635 40103
rect 40785 40069 40819 40103
rect 46857 40069 46891 40103
rect 49249 40069 49283 40103
rect 51273 40069 51307 40103
rect 54033 40069 54067 40103
rect 22477 40001 22511 40035
rect 23581 40001 23615 40035
rect 24665 40001 24699 40035
rect 26249 40001 26283 40035
rect 26433 40001 26467 40035
rect 27905 40001 27939 40035
rect 28181 40001 28215 40035
rect 30665 40001 30699 40035
rect 30849 40001 30883 40035
rect 31033 40001 31067 40035
rect 32873 40001 32907 40035
rect 33021 40001 33055 40035
rect 33338 40001 33372 40035
rect 34713 40001 34747 40035
rect 37749 40001 37783 40035
rect 38393 40001 38427 40035
rect 38577 40001 38611 40035
rect 39681 40001 39715 40035
rect 39773 40001 39807 40035
rect 41521 40001 41555 40035
rect 41705 40001 41739 40035
rect 44097 40001 44131 40035
rect 45109 40001 45143 40035
rect 48053 40001 48087 40035
rect 49893 40001 49927 40035
rect 50077 40001 50111 40035
rect 50629 40001 50663 40035
rect 50813 40001 50847 40035
rect 51549 40001 51583 40035
rect 52929 40001 52963 40035
rect 53941 40001 53975 40035
rect 54125 40001 54159 40035
rect 54769 40001 54803 40035
rect 56149 40001 56183 40035
rect 57897 40001 57931 40035
rect 23673 39933 23707 39967
rect 24409 39933 24443 39967
rect 26341 39933 26375 39967
rect 34897 39933 34931 39967
rect 34989 39933 35023 39967
rect 37565 39933 37599 39967
rect 45201 39933 45235 39967
rect 48237 39933 48271 39967
rect 53021 39933 53055 39967
rect 54861 39933 54895 39967
rect 55137 39933 55171 39967
rect 56241 39933 56275 39967
rect 28917 39865 28951 39899
rect 50721 39865 50755 39899
rect 51825 39865 51859 39899
rect 58081 39865 58115 39899
rect 2421 39797 2455 39831
rect 32321 39797 32355 39831
rect 33517 39797 33551 39831
rect 34529 39797 34563 39831
rect 39497 39797 39531 39831
rect 41521 39797 41555 39831
rect 44281 39797 44315 39831
rect 45385 39797 45419 39831
rect 46949 39797 46983 39831
rect 49341 39797 49375 39831
rect 49985 39797 50019 39831
rect 53205 39797 53239 39831
rect 22845 39593 22879 39627
rect 24409 39593 24443 39627
rect 25697 39593 25731 39627
rect 39865 39593 39899 39627
rect 40325 39593 40359 39627
rect 48421 39593 48455 39627
rect 55781 39593 55815 39627
rect 56425 39593 56459 39627
rect 56793 39593 56827 39627
rect 29009 39525 29043 39559
rect 54769 39525 54803 39559
rect 55597 39525 55631 39559
rect 23857 39457 23891 39491
rect 35173 39457 35207 39491
rect 39957 39457 39991 39491
rect 41061 39457 41095 39491
rect 44465 39457 44499 39491
rect 48881 39457 48915 39491
rect 51181 39457 51215 39491
rect 54493 39457 54527 39491
rect 3801 39389 3835 39423
rect 20913 39389 20947 39423
rect 21097 39389 21131 39423
rect 22753 39389 22787 39423
rect 22937 39389 22971 39423
rect 24639 39389 24673 39423
rect 24777 39389 24811 39423
rect 24874 39389 24908 39423
rect 25053 39389 25087 39423
rect 25605 39389 25639 39423
rect 27629 39389 27663 39423
rect 27896 39389 27930 39423
rect 29929 39389 29963 39423
rect 30757 39389 30791 39423
rect 31769 39389 31803 39423
rect 31917 39389 31951 39423
rect 32137 39389 32171 39423
rect 32275 39389 32309 39423
rect 32873 39389 32907 39423
rect 33021 39389 33055 39423
rect 33149 39389 33183 39423
rect 33357 39389 33391 39423
rect 34897 39389 34931 39423
rect 34989 39389 35023 39423
rect 35081 39389 35115 39423
rect 40141 39389 40175 39423
rect 44281 39389 44315 39423
rect 45293 39389 45327 39423
rect 45385 39389 45419 39423
rect 45477 39389 45511 39423
rect 45661 39389 45695 39423
rect 48605 39389 48639 39423
rect 48697 39389 48731 39423
rect 48973 39389 49007 39423
rect 50169 39389 50203 39423
rect 50905 39389 50939 39423
rect 54401 39389 54435 39423
rect 55321 39389 55355 39423
rect 56333 39389 56367 39423
rect 57253 39389 57287 39423
rect 23673 39321 23707 39355
rect 30849 39321 30883 39355
rect 32045 39321 32079 39355
rect 33241 39321 33275 39355
rect 39865 39321 39899 39355
rect 40877 39321 40911 39355
rect 44097 39321 44131 39355
rect 3893 39253 3927 39287
rect 21097 39253 21131 39287
rect 30021 39253 30055 39287
rect 32413 39253 32447 39287
rect 33517 39253 33551 39287
rect 34713 39253 34747 39287
rect 45017 39253 45051 39287
rect 50353 39253 50387 39287
rect 57345 39253 57379 39287
rect 29009 39049 29043 39083
rect 30773 39049 30807 39083
rect 31493 39049 31527 39083
rect 33057 39049 33091 39083
rect 34345 39049 34379 39083
rect 40969 39049 41003 39083
rect 43453 39049 43487 39083
rect 50169 39049 50203 39083
rect 50951 39049 50985 39083
rect 52101 39049 52135 39083
rect 53481 39049 53515 39083
rect 2421 38981 2455 39015
rect 30573 38981 30607 39015
rect 32689 38981 32723 39015
rect 32781 38981 32815 39015
rect 37565 38981 37599 39015
rect 41705 38981 41739 39015
rect 48513 38981 48547 39015
rect 49985 38981 50019 39015
rect 2237 38913 2271 38947
rect 20913 38913 20947 38947
rect 21005 38913 21039 38947
rect 21097 38913 21131 38947
rect 21281 38913 21315 38947
rect 22017 38913 22051 38947
rect 22753 38913 22787 38947
rect 23857 38913 23891 38947
rect 27997 38913 28031 38947
rect 28273 38913 28307 38947
rect 29469 38913 29503 38947
rect 29653 38913 29687 38947
rect 29929 38913 29963 38947
rect 30113 38913 30147 38947
rect 31401 38913 31435 38947
rect 31585 38913 31619 38947
rect 32413 38913 32447 38947
rect 32506 38913 32540 38947
rect 32919 38913 32953 38947
rect 33517 38913 33551 38947
rect 34529 38913 34563 38947
rect 35357 38913 35391 38947
rect 35541 38913 35575 38947
rect 37289 38913 37323 38947
rect 37473 38913 37507 38947
rect 37657 38913 37691 38947
rect 38393 38913 38427 38947
rect 38577 38913 38611 38947
rect 39776 38913 39810 38947
rect 39865 38913 39899 38947
rect 40049 38913 40083 38947
rect 40151 38913 40185 38947
rect 40601 38913 40635 38947
rect 41521 38913 41555 38947
rect 43637 38913 43671 38947
rect 43729 38913 43763 38947
rect 43913 38913 43947 38947
rect 44005 38913 44039 38947
rect 44741 38913 44775 38947
rect 45017 38913 45051 38947
rect 45201 38913 45235 38947
rect 45937 38913 45971 38947
rect 46029 38913 46063 38947
rect 46121 38913 46155 38947
rect 46305 38913 46339 38947
rect 46857 38913 46891 38947
rect 48329 38913 48363 38947
rect 49341 38913 49375 38947
rect 50261 38913 50295 38947
rect 52009 38913 52043 38947
rect 52193 38913 52227 38947
rect 53297 38913 53331 38947
rect 2789 38845 2823 38879
rect 22293 38845 22327 38879
rect 23029 38845 23063 38879
rect 24593 38845 24627 38879
rect 24869 38845 24903 38879
rect 34621 38845 34655 38879
rect 34713 38845 34747 38879
rect 34805 38845 34839 38879
rect 40693 38845 40727 38879
rect 49433 38845 49467 38879
rect 50721 38845 50755 38879
rect 53113 38845 53147 38879
rect 22845 38777 22879 38811
rect 33609 38777 33643 38811
rect 39589 38777 39623 38811
rect 44833 38777 44867 38811
rect 49985 38777 50019 38811
rect 20637 38709 20671 38743
rect 21833 38709 21867 38743
rect 22201 38709 22235 38743
rect 22937 38709 22971 38743
rect 23949 38709 23983 38743
rect 30757 38709 30791 38743
rect 30941 38709 30975 38743
rect 35357 38709 35391 38743
rect 37841 38709 37875 38743
rect 40601 38709 40635 38743
rect 44465 38709 44499 38743
rect 44925 38709 44959 38743
rect 45661 38709 45695 38743
rect 46949 38709 46983 38743
rect 58081 38709 58115 38743
rect 29561 38505 29595 38539
rect 35725 38505 35759 38539
rect 38485 38505 38519 38539
rect 46305 38505 46339 38539
rect 49525 38505 49559 38539
rect 51641 38505 51675 38539
rect 52653 38505 52687 38539
rect 53021 38505 53055 38539
rect 53665 38505 53699 38539
rect 26709 38437 26743 38471
rect 53573 38437 53607 38471
rect 22753 38369 22787 38403
rect 24869 38369 24903 38403
rect 24961 38369 24995 38403
rect 32413 38369 32447 38403
rect 34989 38369 35023 38403
rect 35173 38369 35207 38403
rect 38761 38369 38795 38403
rect 38853 38369 38887 38403
rect 38945 38369 38979 38403
rect 40417 38369 40451 38403
rect 41337 38369 41371 38403
rect 43913 38369 43947 38403
rect 45293 38369 45327 38403
rect 50169 38369 50203 38403
rect 53757 38369 53791 38403
rect 56333 38369 56367 38403
rect 57897 38369 57931 38403
rect 19257 38301 19291 38335
rect 21925 38301 21959 38335
rect 22017 38301 22051 38335
rect 22130 38298 22164 38332
rect 22293 38301 22327 38335
rect 22937 38301 22971 38335
rect 23213 38301 23247 38335
rect 24777 38301 24811 38335
rect 25053 38301 25087 38335
rect 29745 38301 29779 38335
rect 30021 38301 30055 38335
rect 30205 38301 30239 38335
rect 30665 38301 30699 38335
rect 31033 38301 31067 38335
rect 32689 38301 32723 38335
rect 33701 38301 33735 38335
rect 33885 38301 33919 38335
rect 34897 38301 34931 38335
rect 35081 38301 35115 38335
rect 35725 38301 35759 38335
rect 35909 38301 35943 38335
rect 36461 38301 36495 38335
rect 36645 38301 36679 38335
rect 36829 38301 36863 38335
rect 37473 38301 37507 38335
rect 37841 38301 37875 38335
rect 38669 38301 38703 38335
rect 39865 38301 39899 38335
rect 40325 38301 40359 38335
rect 40693 38301 40727 38335
rect 40785 38301 40819 38335
rect 41521 38301 41555 38335
rect 41797 38301 41831 38335
rect 43269 38301 43303 38335
rect 43453 38301 43487 38335
rect 43637 38301 43671 38335
rect 45017 38301 45051 38335
rect 46581 38301 46615 38335
rect 46670 38295 46704 38329
rect 46770 38301 46804 38335
rect 46949 38301 46983 38335
rect 48329 38301 48363 38335
rect 48513 38301 48547 38335
rect 49433 38301 49467 38335
rect 49617 38301 49651 38335
rect 50445 38301 50479 38335
rect 52653 38301 52687 38335
rect 52837 38301 52871 38335
rect 53481 38301 53515 38335
rect 19524 38233 19558 38267
rect 23121 38233 23155 38267
rect 26525 38233 26559 38267
rect 30849 38233 30883 38267
rect 31585 38233 31619 38267
rect 33793 38233 33827 38267
rect 36737 38233 36771 38267
rect 37657 38233 37691 38267
rect 37749 38233 37783 38267
rect 40049 38233 40083 38267
rect 43545 38233 43579 38267
rect 43755 38233 43789 38267
rect 47501 38233 47535 38267
rect 51457 38233 51491 38267
rect 51657 38233 51691 38267
rect 56517 38233 56551 38267
rect 20637 38165 20671 38199
rect 21649 38165 21683 38199
rect 24593 38165 24627 38199
rect 31677 38165 31711 38199
rect 34713 38165 34747 38199
rect 37013 38165 37047 38199
rect 38025 38165 38059 38199
rect 41705 38165 41739 38199
rect 47593 38165 47627 38199
rect 48421 38165 48455 38199
rect 51825 38165 51859 38199
rect 22017 37961 22051 37995
rect 22661 37961 22695 37995
rect 23121 37961 23155 37995
rect 24593 37961 24627 37995
rect 24685 37961 24719 37995
rect 24869 37961 24903 37995
rect 25529 37961 25563 37995
rect 29653 37961 29687 37995
rect 39957 37961 39991 37995
rect 41245 37961 41279 37995
rect 42533 37961 42567 37995
rect 44005 37961 44039 37995
rect 45753 37961 45787 37995
rect 48973 37961 49007 37995
rect 52193 37961 52227 37995
rect 25329 37893 25363 37927
rect 36369 37893 36403 37927
rect 43637 37893 43671 37927
rect 44465 37893 44499 37927
rect 47777 37893 47811 37927
rect 51825 37893 51859 37927
rect 52025 37893 52059 37927
rect 20085 37825 20119 37859
rect 21005 37825 21039 37859
rect 22477 37825 22511 37859
rect 23581 37825 23615 37859
rect 24501 37825 24535 37859
rect 24869 37825 24903 37859
rect 26341 37825 26375 37859
rect 29929 37825 29963 37859
rect 30757 37825 30791 37859
rect 32505 37825 32539 37859
rect 33517 37825 33551 37859
rect 34805 37825 34839 37859
rect 36205 37825 36239 37859
rect 36461 37825 36495 37859
rect 36553 37825 36587 37859
rect 37565 37825 37599 37859
rect 38577 37825 38611 37859
rect 38761 37825 38795 37859
rect 38853 37825 38887 37859
rect 38945 37825 38979 37859
rect 40141 37825 40175 37859
rect 40233 37825 40267 37859
rect 40509 37825 40543 37859
rect 41429 37825 41463 37859
rect 41521 37825 41555 37859
rect 41797 37825 41831 37859
rect 42441 37825 42475 37859
rect 42717 37825 42751 37859
rect 43810 37825 43844 37859
rect 44649 37825 44683 37859
rect 46305 37825 46339 37859
rect 46489 37825 46523 37859
rect 47593 37825 47627 37859
rect 48789 37825 48823 37859
rect 48881 37825 48915 37859
rect 49801 37825 49835 37859
rect 49985 37825 50019 37859
rect 50077 37825 50111 37859
rect 50813 37825 50847 37859
rect 53113 37825 53147 37859
rect 56793 37825 56827 37859
rect 20177 37757 20211 37791
rect 22385 37757 22419 37791
rect 23305 37757 23339 37791
rect 23397 37757 23431 37791
rect 23489 37757 23523 37791
rect 29837 37757 29871 37791
rect 30021 37757 30055 37791
rect 30113 37757 30147 37791
rect 31033 37757 31067 37791
rect 32413 37757 32447 37791
rect 32597 37757 32631 37791
rect 32689 37757 32723 37791
rect 33241 37757 33275 37791
rect 34529 37757 34563 37791
rect 37289 37757 37323 37791
rect 41705 37757 41739 37791
rect 44833 37757 44867 37791
rect 44925 37757 44959 37791
rect 46029 37757 46063 37791
rect 50537 37757 50571 37791
rect 53205 37757 53239 37791
rect 56885 37757 56919 37791
rect 57161 37757 57195 37791
rect 25697 37689 25731 37723
rect 46121 37689 46155 37723
rect 48605 37689 48639 37723
rect 49157 37689 49191 37723
rect 53481 37689 53515 37723
rect 20453 37621 20487 37655
rect 21189 37621 21223 37655
rect 25513 37621 25547 37655
rect 26157 37621 26191 37655
rect 32229 37621 32263 37655
rect 36737 37621 36771 37655
rect 39129 37621 39163 37655
rect 40417 37621 40451 37655
rect 46213 37621 46247 37655
rect 47961 37621 47995 37655
rect 49801 37621 49835 37655
rect 52009 37621 52043 37655
rect 20637 37417 20671 37451
rect 23397 37417 23431 37451
rect 28273 37417 28307 37451
rect 30297 37417 30331 37451
rect 42993 37417 43027 37451
rect 45385 37417 45419 37451
rect 45937 37417 45971 37451
rect 47225 37417 47259 37451
rect 47409 37417 47443 37451
rect 47869 37417 47903 37451
rect 40141 37349 40175 37383
rect 57805 37349 57839 37383
rect 20453 37281 20487 37315
rect 31677 37281 31711 37315
rect 33333 37281 33367 37315
rect 34989 37281 35023 37315
rect 36553 37281 36587 37315
rect 36829 37281 36863 37315
rect 43637 37281 43671 37315
rect 45477 37281 45511 37315
rect 50353 37281 50387 37315
rect 50537 37281 50571 37315
rect 56609 37281 56643 37315
rect 57253 37281 57287 37315
rect 20361 37213 20395 37247
rect 21373 37213 21407 37247
rect 23213 37213 23247 37247
rect 25881 37213 25915 37247
rect 28181 37213 28215 37247
rect 30481 37213 30515 37247
rect 30573 37213 30607 37247
rect 31401 37213 31435 37247
rect 31585 37213 31619 37247
rect 31815 37213 31849 37247
rect 31953 37213 31987 37247
rect 33609 37213 33643 37247
rect 34713 37213 34747 37247
rect 37841 37213 37875 37247
rect 38209 37213 38243 37247
rect 40601 37213 40635 37247
rect 40969 37213 41003 37247
rect 45201 37213 45235 37247
rect 45937 37213 45971 37247
rect 46121 37213 46155 37247
rect 46213 37213 46247 37247
rect 48145 37213 48179 37247
rect 48881 37213 48915 37247
rect 49157 37213 49191 37247
rect 49249 37213 49283 37247
rect 50445 37213 50479 37247
rect 50629 37213 50663 37247
rect 56701 37213 56735 37247
rect 58081 37213 58115 37247
rect 21640 37145 21674 37179
rect 26148 37145 26182 37179
rect 30297 37145 30331 37179
rect 38025 37145 38059 37179
rect 38117 37145 38151 37179
rect 39957 37145 39991 37179
rect 40785 37145 40819 37179
rect 40877 37145 40911 37179
rect 43361 37145 43395 37179
rect 47041 37145 47075 37179
rect 47257 37145 47291 37179
rect 47869 37145 47903 37179
rect 49065 37145 49099 37179
rect 57805 37145 57839 37179
rect 22753 37077 22787 37111
rect 27261 37077 27295 37111
rect 32137 37077 32171 37111
rect 38393 37077 38427 37111
rect 41153 37077 41187 37111
rect 43453 37077 43487 37111
rect 45017 37077 45051 37111
rect 48053 37077 48087 37111
rect 49433 37077 49467 37111
rect 50169 37077 50203 37111
rect 57989 37077 58023 37111
rect 23121 36873 23155 36907
rect 33517 36873 33551 36907
rect 44833 36873 44867 36907
rect 49065 36873 49099 36907
rect 50169 36873 50203 36907
rect 56425 36873 56459 36907
rect 57345 36873 57379 36907
rect 57989 36873 58023 36907
rect 31125 36805 31159 36839
rect 36369 36805 36403 36839
rect 37473 36805 37507 36839
rect 37565 36805 37599 36839
rect 48605 36805 48639 36839
rect 49801 36805 49835 36839
rect 50031 36771 50065 36805
rect 22017 36737 22051 36771
rect 22845 36737 22879 36771
rect 22937 36737 22971 36771
rect 25973 36737 26007 36771
rect 28457 36737 28491 36771
rect 29377 36737 29411 36771
rect 33425 36737 33459 36771
rect 33609 36737 33643 36771
rect 34253 36737 34287 36771
rect 34529 36737 34563 36771
rect 35265 36737 35299 36771
rect 36185 36737 36219 36771
rect 36461 36737 36495 36771
rect 36553 36737 36587 36771
rect 37289 36737 37323 36771
rect 37657 36737 37691 36771
rect 40969 36737 41003 36771
rect 44465 36737 44499 36771
rect 44557 36737 44591 36771
rect 47777 36737 47811 36771
rect 48881 36737 48915 36771
rect 50629 36737 50663 36771
rect 50813 36737 50847 36771
rect 54033 36737 54067 36771
rect 55045 36737 55079 36771
rect 56057 36737 56091 36771
rect 56885 36737 56919 36771
rect 57897 36737 57931 36771
rect 22109 36669 22143 36703
rect 23121 36669 23155 36703
rect 26249 36669 26283 36703
rect 28733 36669 28767 36703
rect 29193 36669 29227 36703
rect 29653 36669 29687 36703
rect 34345 36669 34379 36703
rect 34437 36669 34471 36703
rect 35357 36669 35391 36703
rect 35449 36669 35483 36703
rect 35541 36669 35575 36703
rect 47593 36669 47627 36703
rect 48697 36669 48731 36703
rect 53941 36669 53975 36703
rect 54953 36669 54987 36703
rect 55965 36669 55999 36703
rect 22385 36601 22419 36635
rect 31309 36601 31343 36635
rect 41153 36601 41187 36635
rect 54401 36601 54435 36635
rect 55413 36601 55447 36635
rect 25789 36533 25823 36567
rect 26157 36533 26191 36567
rect 28273 36533 28307 36567
rect 28641 36533 28675 36567
rect 29561 36533 29595 36567
rect 34069 36533 34103 36567
rect 35081 36533 35115 36567
rect 36737 36533 36771 36567
rect 37841 36533 37875 36567
rect 44649 36533 44683 36567
rect 47961 36533 47995 36567
rect 48881 36533 48915 36567
rect 49985 36533 50019 36567
rect 50629 36533 50663 36567
rect 57161 36533 57195 36567
rect 26617 36329 26651 36363
rect 33977 36329 34011 36363
rect 35725 36329 35759 36363
rect 43453 36329 43487 36363
rect 45569 36329 45603 36363
rect 46029 36329 46063 36363
rect 47593 36329 47627 36363
rect 53665 36329 53699 36363
rect 56425 36329 56459 36363
rect 57253 36329 57287 36363
rect 44005 36261 44039 36295
rect 46857 36261 46891 36295
rect 48329 36261 48363 36295
rect 52745 36261 52779 36295
rect 29561 36193 29595 36227
rect 29837 36193 29871 36227
rect 33057 36193 33091 36227
rect 34897 36193 34931 36227
rect 35081 36193 35115 36227
rect 43269 36193 43303 36227
rect 45937 36193 45971 36227
rect 48053 36193 48087 36227
rect 52285 36193 52319 36227
rect 53297 36193 53331 36227
rect 56149 36193 56183 36227
rect 24409 36125 24443 36159
rect 26433 36125 26467 36159
rect 26709 36125 26743 36159
rect 27537 36125 27571 36159
rect 27804 36125 27838 36159
rect 30941 36125 30975 36159
rect 32873 36125 32907 36159
rect 33977 36125 34011 36159
rect 34161 36125 34195 36159
rect 34989 36125 35023 36159
rect 35173 36125 35207 36159
rect 35725 36125 35759 36159
rect 35909 36125 35943 36159
rect 43177 36125 43211 36159
rect 44281 36125 44315 36159
rect 45845 36125 45879 36159
rect 46121 36125 46155 36159
rect 46305 36125 46339 36159
rect 48237 36125 48271 36159
rect 48605 36125 48639 36159
rect 52377 36125 52411 36159
rect 53389 36125 53423 36159
rect 56057 36125 56091 36159
rect 56885 36125 56919 36159
rect 24676 36057 24710 36091
rect 31208 36057 31242 36091
rect 44005 36057 44039 36091
rect 46857 36057 46891 36091
rect 47317 36057 47351 36091
rect 57069 36057 57103 36091
rect 25789 35989 25823 36023
rect 26249 35989 26283 36023
rect 28917 35989 28951 36023
rect 32321 35989 32355 36023
rect 34713 35989 34747 36023
rect 44189 35989 44223 36023
rect 47409 35989 47443 36023
rect 48513 35989 48547 36023
rect 26985 35785 27019 35819
rect 32689 35785 32723 35819
rect 43821 35785 43855 35819
rect 48145 35785 48179 35819
rect 25320 35717 25354 35751
rect 31309 35717 31343 35751
rect 32597 35717 32631 35751
rect 43453 35717 43487 35751
rect 45293 35717 45327 35751
rect 49801 35717 49835 35751
rect 50001 35717 50035 35751
rect 51641 35717 51675 35751
rect 55229 35717 55263 35751
rect 25053 35649 25087 35683
rect 27169 35649 27203 35683
rect 27905 35649 27939 35683
rect 28172 35649 28206 35683
rect 31217 35649 31251 35683
rect 34345 35649 34379 35683
rect 34437 35649 34471 35683
rect 35173 35649 35207 35683
rect 35357 35649 35391 35683
rect 37545 35649 37579 35683
rect 40417 35649 40451 35683
rect 41429 35649 41463 35683
rect 42809 35649 42843 35683
rect 42993 35649 43027 35683
rect 43637 35649 43671 35683
rect 44281 35649 44315 35683
rect 44465 35649 44499 35683
rect 45109 35649 45143 35683
rect 45385 35649 45419 35683
rect 48053 35649 48087 35683
rect 50721 35649 50755 35683
rect 51457 35649 51491 35683
rect 51733 35649 51767 35683
rect 55413 35649 55447 35683
rect 56149 35649 56183 35683
rect 27445 35581 27479 35615
rect 31493 35581 31527 35615
rect 34529 35581 34563 35615
rect 34621 35581 34655 35615
rect 37289 35581 37323 35615
rect 40509 35581 40543 35615
rect 41705 35581 41739 35615
rect 27353 35513 27387 35547
rect 41245 35513 41279 35547
rect 26433 35445 26467 35479
rect 29285 35445 29319 35479
rect 30849 35445 30883 35479
rect 34161 35445 34195 35479
rect 35173 35445 35207 35479
rect 38669 35445 38703 35479
rect 40693 35445 40727 35479
rect 41613 35445 41647 35479
rect 42901 35445 42935 35479
rect 44649 35445 44683 35479
rect 45109 35445 45143 35479
rect 49985 35445 50019 35479
rect 50169 35445 50203 35479
rect 50813 35445 50847 35479
rect 51457 35445 51491 35479
rect 55597 35445 55631 35479
rect 56241 35445 56275 35479
rect 56609 35445 56643 35479
rect 27353 35241 27387 35275
rect 32413 35241 32447 35275
rect 40509 35241 40543 35275
rect 41889 35241 41923 35275
rect 47225 35241 47259 35275
rect 49249 35241 49283 35275
rect 50721 35241 50755 35275
rect 52193 35241 52227 35275
rect 57253 35241 57287 35275
rect 26249 35173 26283 35207
rect 29837 35173 29871 35207
rect 46121 35173 46155 35207
rect 24869 35105 24903 35139
rect 28181 35105 28215 35139
rect 30481 35105 30515 35139
rect 31033 35105 31067 35139
rect 34713 35105 34747 35139
rect 40969 35105 41003 35139
rect 41061 35105 41095 35139
rect 43085 35105 43119 35139
rect 43637 35105 43671 35139
rect 43729 35105 43763 35139
rect 44373 35105 44407 35139
rect 51273 35105 51307 35139
rect 52561 35105 52595 35139
rect 25136 35037 25170 35071
rect 27261 35037 27295 35071
rect 28457 35037 28491 35071
rect 30297 35037 30331 35071
rect 37197 35037 37231 35071
rect 37464 35037 37498 35071
rect 41705 35037 41739 35071
rect 42717 35037 42751 35071
rect 42993 35037 43027 35071
rect 44097 35037 44131 35071
rect 45661 35037 45695 35071
rect 46397 35037 46431 35071
rect 47133 35037 47167 35071
rect 47317 35037 47351 35071
rect 51089 35037 51123 35071
rect 52377 35037 52411 35071
rect 52469 35037 52503 35071
rect 52653 35037 52687 35071
rect 53205 35037 53239 35071
rect 53389 35037 53423 35071
rect 56241 35037 56275 35071
rect 56425 35037 56459 35071
rect 56977 35037 57011 35071
rect 57069 35037 57103 35071
rect 31300 34969 31334 35003
rect 34980 34969 35014 35003
rect 40877 34969 40911 35003
rect 44189 34969 44223 35003
rect 45477 34969 45511 35003
rect 46121 34969 46155 35003
rect 49157 34969 49191 35003
rect 30205 34901 30239 34935
rect 36093 34901 36127 34935
rect 38577 34901 38611 34935
rect 46305 34901 46339 34935
rect 51181 34901 51215 34935
rect 53297 34901 53331 34935
rect 56425 34901 56459 34935
rect 31585 34697 31619 34731
rect 38669 34697 38703 34731
rect 41061 34697 41095 34731
rect 42993 34697 43027 34731
rect 43361 34697 43395 34731
rect 44373 34697 44407 34731
rect 46489 34697 46523 34731
rect 49065 34697 49099 34731
rect 51917 34697 51951 34731
rect 52929 34697 52963 34731
rect 37556 34629 37590 34663
rect 41705 34629 41739 34663
rect 43913 34629 43947 34663
rect 45937 34629 45971 34663
rect 49801 34629 49835 34663
rect 50077 34629 50111 34663
rect 50721 34629 50755 34663
rect 50813 34629 50847 34663
rect 28181 34561 28215 34595
rect 30205 34561 30239 34595
rect 30472 34561 30506 34595
rect 32321 34561 32355 34595
rect 32597 34561 32631 34595
rect 33241 34561 33275 34595
rect 34069 34561 34103 34595
rect 34325 34561 34359 34595
rect 37289 34561 37323 34595
rect 40417 34561 40451 34595
rect 40693 34561 40727 34595
rect 41521 34561 41555 34595
rect 43177 34561 43211 34595
rect 43453 34561 43487 34595
rect 44189 34561 44223 34595
rect 44925 34561 44959 34595
rect 45201 34561 45235 34595
rect 45845 34561 45879 34595
rect 46029 34561 46063 34595
rect 46673 34561 46707 34595
rect 46857 34561 46891 34595
rect 47869 34561 47903 34595
rect 48881 34561 48915 34595
rect 49065 34561 49099 34595
rect 49525 34561 49559 34595
rect 49709 34561 49743 34595
rect 49893 34561 49927 34595
rect 50537 34561 50571 34595
rect 50905 34561 50939 34595
rect 51733 34561 51767 34595
rect 52009 34561 52043 34595
rect 52745 34561 52779 34595
rect 56885 34561 56919 34595
rect 27997 34493 28031 34527
rect 32505 34493 32539 34527
rect 44097 34493 44131 34527
rect 45017 34493 45051 34527
rect 46765 34493 46799 34527
rect 46949 34493 46983 34527
rect 47593 34493 47627 34527
rect 51549 34493 51583 34527
rect 32137 34425 32171 34459
rect 35449 34425 35483 34459
rect 28365 34357 28399 34391
rect 33057 34357 33091 34391
rect 41889 34357 41923 34391
rect 44189 34357 44223 34391
rect 44925 34357 44959 34391
rect 45385 34357 45419 34391
rect 51089 34357 51123 34391
rect 56977 34357 57011 34391
rect 58081 34357 58115 34391
rect 28181 34153 28215 34187
rect 39129 34153 39163 34187
rect 40325 34153 40359 34187
rect 44097 34153 44131 34187
rect 45201 34153 45235 34187
rect 47225 34153 47259 34187
rect 51273 34153 51307 34187
rect 52009 34153 52043 34187
rect 52193 34153 52227 34187
rect 54493 34153 54527 34187
rect 55873 34153 55907 34187
rect 43729 34085 43763 34119
rect 44281 34085 44315 34119
rect 45385 34085 45419 34119
rect 25513 34017 25547 34051
rect 25697 34017 25731 34051
rect 28641 34017 28675 34051
rect 28825 34017 28859 34051
rect 30757 34017 30791 34051
rect 34713 34017 34747 34051
rect 39037 34017 39071 34051
rect 40969 34017 41003 34051
rect 41521 34017 41555 34051
rect 41981 34017 42015 34051
rect 44189 34017 44223 34051
rect 47501 34017 47535 34051
rect 47685 34017 47719 34051
rect 53481 34017 53515 34051
rect 56333 34017 56367 34051
rect 56517 34017 56551 34051
rect 57897 34017 57931 34051
rect 27721 33949 27755 33983
rect 34969 33949 35003 33983
rect 38945 33949 38979 33983
rect 41889 33949 41923 33983
rect 44005 33949 44039 33983
rect 44465 33949 44499 33983
rect 46489 33949 46523 33983
rect 46765 33949 46799 33983
rect 47409 33949 47443 33983
rect 47593 33949 47627 33983
rect 48421 33949 48455 33983
rect 52653 33949 52687 33983
rect 52837 33949 52871 33983
rect 53573 33949 53607 33983
rect 54493 33949 54527 33983
rect 54677 33949 54711 33983
rect 55597 33949 55631 33983
rect 55689 33949 55723 33983
rect 25421 33881 25455 33915
rect 31002 33881 31036 33915
rect 40785 33881 40819 33915
rect 42165 33881 42199 33915
rect 42717 33881 42751 33915
rect 45017 33881 45051 33915
rect 45233 33881 45267 33915
rect 46305 33881 46339 33915
rect 49341 33881 49375 33915
rect 49525 33881 49559 33915
rect 50997 33881 51031 33915
rect 51825 33881 51859 33915
rect 52745 33881 52779 33915
rect 25053 33813 25087 33847
rect 27537 33813 27571 33847
rect 28549 33813 28583 33847
rect 32137 33813 32171 33847
rect 36093 33813 36127 33847
rect 39313 33813 39347 33847
rect 40693 33813 40727 33847
rect 42809 33813 42843 33847
rect 46673 33813 46707 33847
rect 48513 33813 48547 33847
rect 52025 33813 52059 33847
rect 53941 33813 53975 33847
rect 26065 33609 26099 33643
rect 30757 33609 30791 33643
rect 41613 33609 41647 33643
rect 42993 33609 43027 33643
rect 44281 33609 44315 33643
rect 45569 33609 45603 33643
rect 47685 33609 47719 33643
rect 47869 33609 47903 33643
rect 49893 33609 49927 33643
rect 51549 33609 51583 33643
rect 55045 33609 55079 33643
rect 55873 33609 55907 33643
rect 27782 33541 27816 33575
rect 29929 33541 29963 33575
rect 30113 33541 30147 33575
rect 40969 33541 41003 33575
rect 42625 33541 42659 33575
rect 42717 33541 42751 33575
rect 43913 33541 43947 33575
rect 44129 33541 44163 33575
rect 49801 33541 49835 33575
rect 53941 33541 53975 33575
rect 54157 33541 54191 33575
rect 56333 33541 56367 33575
rect 24133 33473 24167 33507
rect 24777 33473 24811 33507
rect 24961 33473 24995 33507
rect 25973 33473 26007 33507
rect 30941 33473 30975 33507
rect 42441 33473 42475 33507
rect 42809 33473 42843 33507
rect 44741 33473 44775 33507
rect 44925 33473 44959 33507
rect 45017 33473 45051 33507
rect 45477 33473 45511 33507
rect 45661 33473 45695 33507
rect 47593 33473 47627 33507
rect 47961 33473 47995 33507
rect 49065 33473 49099 33507
rect 49249 33473 49283 33507
rect 50629 33473 50663 33507
rect 51365 33473 51399 33507
rect 51549 33473 51583 33507
rect 54769 33473 54803 33507
rect 55505 33473 55539 33507
rect 56517 33473 56551 33507
rect 56609 33473 56643 33507
rect 57069 33473 57103 33507
rect 23949 33405 23983 33439
rect 26157 33405 26191 33439
rect 27537 33405 27571 33439
rect 41337 33405 41371 33439
rect 41429 33405 41463 33439
rect 47777 33405 47811 33439
rect 49157 33405 49191 33439
rect 50813 33405 50847 33439
rect 50905 33405 50939 33439
rect 55045 33405 55079 33439
rect 55597 33405 55631 33439
rect 25605 33337 25639 33371
rect 44741 33337 44775 33371
rect 50445 33337 50479 33371
rect 54309 33337 54343 33371
rect 54861 33337 54895 33371
rect 24317 33269 24351 33303
rect 25145 33269 25179 33303
rect 28917 33269 28951 33303
rect 44097 33269 44131 33303
rect 54125 33269 54159 33303
rect 55505 33269 55539 33303
rect 56333 33269 56367 33303
rect 57161 33269 57195 33303
rect 58081 33269 58115 33303
rect 26249 33065 26283 33099
rect 41337 33065 41371 33099
rect 42717 33065 42751 33099
rect 44097 33065 44131 33099
rect 46581 33065 46615 33099
rect 47133 33065 47167 33099
rect 48237 33065 48271 33099
rect 51089 33065 51123 33099
rect 53849 33065 53883 33099
rect 55689 33065 55723 33099
rect 48421 32997 48455 33031
rect 51273 32997 51307 33031
rect 51733 32997 51767 33031
rect 26709 32929 26743 32963
rect 26893 32929 26927 32963
rect 27629 32929 27663 32963
rect 30021 32929 30055 32963
rect 30113 32929 30147 32963
rect 50445 32929 50479 32963
rect 56333 32929 56367 32963
rect 56517 32929 56551 32963
rect 57805 32929 57839 32963
rect 23857 32861 23891 32895
rect 24409 32861 24443 32895
rect 36829 32861 36863 32895
rect 37096 32861 37130 32895
rect 41521 32861 41555 32895
rect 41613 32861 41647 32895
rect 41797 32861 41831 32895
rect 41889 32861 41923 32895
rect 44097 32861 44131 32895
rect 44281 32861 44315 32895
rect 45477 32861 45511 32895
rect 45661 32861 45695 32895
rect 46489 32861 46523 32895
rect 46673 32861 46707 32895
rect 47317 32861 47351 32895
rect 47593 32861 47627 32895
rect 51917 32861 51951 32895
rect 52009 32861 52043 32895
rect 54125 32861 54159 32895
rect 54585 32861 54619 32895
rect 54769 32861 54803 32895
rect 48283 32827 48317 32861
rect 24654 32793 24688 32827
rect 27896 32793 27930 32827
rect 29929 32793 29963 32827
rect 42349 32793 42383 32827
rect 42533 32793 42567 32827
rect 48053 32793 48087 32827
rect 50261 32793 50295 32827
rect 50905 32793 50939 32827
rect 51105 32793 51139 32827
rect 51733 32793 51767 32827
rect 53849 32793 53883 32827
rect 54677 32793 54711 32827
rect 55505 32793 55539 32827
rect 55721 32793 55755 32827
rect 23673 32725 23707 32759
rect 25789 32725 25823 32759
rect 26617 32725 26651 32759
rect 29009 32725 29043 32759
rect 29561 32725 29595 32759
rect 38209 32725 38243 32759
rect 45569 32725 45603 32759
rect 47501 32725 47535 32759
rect 54033 32725 54067 32759
rect 55873 32725 55907 32759
rect 26249 32521 26283 32555
rect 41061 32521 41095 32555
rect 41429 32521 41463 32555
rect 42441 32521 42475 32555
rect 47685 32521 47719 32555
rect 52745 32521 52779 32555
rect 53573 32521 53607 32555
rect 56517 32521 56551 32555
rect 57069 32521 57103 32555
rect 37534 32453 37568 32487
rect 48697 32453 48731 32487
rect 51089 32453 51123 32487
rect 51825 32453 51859 32487
rect 24041 32385 24075 32419
rect 24225 32385 24259 32419
rect 24869 32385 24903 32419
rect 25136 32385 25170 32419
rect 27169 32385 27203 32419
rect 28825 32385 28859 32419
rect 32321 32385 32355 32419
rect 34161 32385 34195 32419
rect 34428 32385 34462 32419
rect 37289 32385 37323 32419
rect 41245 32385 41279 32419
rect 41521 32385 41555 32419
rect 42625 32385 42659 32419
rect 42717 32385 42751 32419
rect 42901 32385 42935 32419
rect 42993 32385 43027 32419
rect 45017 32385 45051 32419
rect 45201 32385 45235 32419
rect 47869 32385 47903 32419
rect 47961 32385 47995 32419
rect 48145 32385 48179 32419
rect 48237 32385 48271 32419
rect 48881 32385 48915 32419
rect 49985 32385 50019 32419
rect 50169 32385 50203 32419
rect 50905 32385 50939 32419
rect 52009 32385 52043 32419
rect 52745 32385 52779 32419
rect 53481 32385 53515 32419
rect 53665 32385 53699 32419
rect 56241 32385 56275 32419
rect 56977 32385 57011 32419
rect 57161 32385 57195 32419
rect 28641 32317 28675 32351
rect 32137 32317 32171 32351
rect 49065 32317 49099 32351
rect 53021 32317 53055 32351
rect 55873 32317 55907 32351
rect 56333 32317 56367 32351
rect 50077 32249 50111 32283
rect 52837 32249 52871 32283
rect 24409 32181 24443 32215
rect 26985 32181 27019 32215
rect 29009 32181 29043 32215
rect 32505 32181 32539 32215
rect 35541 32181 35575 32215
rect 38669 32181 38703 32215
rect 45109 32181 45143 32215
rect 52193 32181 52227 32215
rect 28549 31977 28583 32011
rect 32965 31977 32999 32011
rect 41797 31977 41831 32011
rect 42901 31977 42935 32011
rect 47041 31977 47075 32011
rect 48881 31977 48915 32011
rect 52285 31977 52319 32011
rect 53573 31977 53607 32011
rect 26433 31909 26467 31943
rect 38577 31909 38611 31943
rect 48145 31909 48179 31943
rect 53205 31909 53239 31943
rect 25053 31841 25087 31875
rect 30297 31841 30331 31875
rect 34713 31841 34747 31875
rect 37197 31841 37231 31875
rect 43545 31841 43579 31875
rect 44373 31841 44407 31875
rect 45293 31841 45327 31875
rect 50629 31841 50663 31875
rect 52745 31841 52779 31875
rect 55689 31841 55723 31875
rect 28733 31773 28767 31807
rect 30481 31773 30515 31807
rect 30665 31773 30699 31807
rect 31125 31773 31159 31807
rect 33149 31773 33183 31807
rect 34969 31773 35003 31807
rect 37464 31773 37498 31807
rect 41981 31773 42015 31807
rect 42165 31773 42199 31807
rect 42257 31773 42291 31807
rect 42809 31773 42843 31807
rect 43453 31773 43487 31807
rect 43637 31773 43671 31807
rect 44281 31773 44315 31807
rect 44465 31773 44499 31807
rect 45477 31773 45511 31807
rect 45661 31773 45695 31807
rect 47225 31773 47259 31807
rect 47409 31773 47443 31807
rect 47501 31773 47535 31807
rect 47961 31773 47995 31807
rect 50905 31773 50939 31807
rect 52469 31773 52503 31807
rect 52653 31773 52687 31807
rect 53389 31773 53423 31807
rect 53665 31773 53699 31807
rect 55873 31773 55907 31807
rect 56057 31773 56091 31807
rect 25320 31705 25354 31739
rect 31370 31705 31404 31739
rect 48789 31705 48823 31739
rect 32505 31637 32539 31671
rect 36093 31637 36127 31671
rect 25053 31433 25087 31467
rect 28733 31433 28767 31467
rect 32137 31433 32171 31467
rect 39865 31433 39899 31467
rect 40509 31433 40543 31467
rect 43269 31433 43303 31467
rect 46673 31433 46707 31467
rect 48145 31433 48179 31467
rect 49709 31433 49743 31467
rect 50997 31433 51031 31467
rect 51365 31433 51399 31467
rect 53481 31433 53515 31467
rect 55597 31433 55631 31467
rect 55965 31433 55999 31467
rect 56609 31433 56643 31467
rect 28825 31365 28859 31399
rect 32597 31365 32631 31399
rect 37556 31365 37590 31399
rect 51181 31365 51215 31399
rect 51825 31365 51859 31399
rect 52929 31365 52963 31399
rect 53757 31365 53791 31399
rect 55045 31365 55079 31399
rect 56701 31365 56735 31399
rect 25237 31297 25271 31331
rect 27537 31297 27571 31331
rect 27721 31297 27755 31331
rect 30389 31297 30423 31331
rect 31217 31297 31251 31331
rect 31309 31297 31343 31331
rect 32505 31297 32539 31331
rect 34989 31297 35023 31331
rect 35256 31297 35290 31331
rect 37289 31297 37323 31331
rect 39497 31297 39531 31331
rect 39681 31297 39715 31331
rect 40417 31297 40451 31331
rect 43453 31297 43487 31331
rect 43729 31297 43763 31331
rect 44189 31297 44223 31331
rect 44373 31297 44407 31331
rect 44833 31297 44867 31331
rect 46121 31297 46155 31331
rect 47593 31297 47627 31331
rect 47961 31297 47995 31331
rect 49157 31297 49191 31331
rect 49341 31297 49375 31331
rect 49433 31297 49467 31331
rect 49525 31297 49559 31331
rect 50169 31297 50203 31331
rect 50353 31297 50387 31331
rect 51089 31297 51123 31331
rect 52009 31297 52043 31331
rect 52101 31297 52135 31331
rect 52745 31297 52779 31331
rect 53021 31297 53055 31331
rect 53481 31297 53515 31331
rect 53573 31297 53607 31331
rect 54953 31297 54987 31331
rect 55137 31297 55171 31331
rect 55781 31297 55815 31331
rect 56057 31297 56091 31331
rect 56517 31297 56551 31331
rect 56793 31297 56827 31331
rect 28917 31229 28951 31263
rect 31401 31229 31435 31263
rect 32689 31229 32723 31263
rect 45109 31229 45143 31263
rect 46397 31229 46431 31263
rect 50261 31229 50295 31263
rect 38669 31161 38703 31195
rect 43637 31161 43671 31195
rect 50813 31161 50847 31195
rect 51825 31161 51859 31195
rect 52745 31161 52779 31195
rect 27905 31093 27939 31127
rect 28365 31093 28399 31127
rect 30205 31093 30239 31127
rect 30849 31093 30883 31127
rect 36369 31093 36403 31127
rect 39497 31093 39531 31127
rect 44189 31093 44223 31127
rect 46489 31093 46523 31127
rect 47961 31093 47995 31127
rect 58081 31093 58115 31127
rect 28273 30889 28307 30923
rect 32413 30889 32447 30923
rect 36737 30889 36771 30923
rect 39037 30889 39071 30923
rect 44281 30889 44315 30923
rect 46305 30889 46339 30923
rect 48237 30889 48271 30923
rect 49157 30889 49191 30923
rect 50721 30889 50755 30923
rect 51365 30889 51399 30923
rect 52285 30889 52319 30923
rect 52469 30889 52503 30923
rect 55781 30889 55815 30923
rect 49019 30821 49053 30855
rect 28917 30753 28951 30787
rect 38945 30753 38979 30787
rect 40233 30753 40267 30787
rect 45293 30753 45327 30787
rect 56333 30753 56367 30787
rect 27721 30685 27755 30719
rect 28733 30685 28767 30719
rect 31033 30685 31067 30719
rect 35725 30685 35759 30719
rect 36645 30685 36679 30719
rect 37565 30685 37599 30719
rect 38853 30685 38887 30719
rect 39129 30685 39163 30719
rect 39957 30685 39991 30719
rect 41245 30685 41279 30719
rect 43453 30685 43487 30719
rect 43637 30685 43671 30719
rect 44097 30685 44131 30719
rect 44281 30685 44315 30719
rect 45017 30685 45051 30719
rect 46489 30685 46523 30719
rect 46765 30685 46799 30719
rect 48145 30685 48179 30719
rect 48881 30685 48915 30719
rect 49341 30685 49375 30719
rect 51273 30685 51307 30719
rect 51457 30685 51491 30719
rect 54493 30685 54527 30719
rect 54677 30685 54711 30719
rect 55597 30685 55631 30719
rect 31278 30617 31312 30651
rect 36001 30617 36035 30651
rect 50629 30617 50663 30651
rect 52101 30617 52135 30651
rect 52317 30617 52351 30651
rect 55413 30617 55447 30651
rect 56517 30617 56551 30651
rect 58173 30617 58207 30651
rect 27537 30549 27571 30583
rect 28641 30549 28675 30583
rect 37105 30549 37139 30583
rect 37749 30549 37783 30583
rect 39313 30549 39347 30583
rect 41337 30549 41371 30583
rect 43545 30549 43579 30583
rect 44465 30549 44499 30583
rect 46673 30549 46707 30583
rect 49341 30549 49375 30583
rect 54585 30549 54619 30583
rect 28365 30345 28399 30379
rect 38669 30345 38703 30379
rect 40325 30345 40359 30379
rect 49525 30345 49559 30379
rect 55781 30345 55815 30379
rect 27252 30277 27286 30311
rect 34152 30277 34186 30311
rect 36645 30277 36679 30311
rect 41889 30277 41923 30311
rect 43269 30277 43303 30311
rect 44373 30277 44407 30311
rect 44833 30277 44867 30311
rect 48973 30277 49007 30311
rect 55597 30277 55631 30311
rect 57989 30277 58023 30311
rect 2421 30209 2455 30243
rect 25973 30209 26007 30243
rect 26985 30209 27019 30243
rect 29009 30209 29043 30243
rect 30849 30209 30883 30243
rect 33885 30209 33919 30243
rect 36461 30209 36495 30243
rect 36737 30209 36771 30243
rect 37565 30209 37599 30243
rect 38393 30209 38427 30243
rect 38853 30209 38887 30243
rect 39313 30209 39347 30243
rect 39957 30209 39991 30243
rect 41521 30209 41555 30243
rect 41705 30209 41739 30243
rect 42441 30209 42475 30243
rect 42533 30209 42567 30243
rect 42809 30209 42843 30243
rect 43453 30209 43487 30243
rect 44189 30209 44223 30243
rect 45017 30209 45051 30243
rect 45201 30209 45235 30243
rect 45293 30209 45327 30243
rect 48053 30209 48087 30243
rect 48237 30209 48271 30243
rect 48789 30209 48823 30243
rect 49433 30209 49467 30243
rect 49617 30209 49651 30243
rect 51089 30209 51123 30243
rect 54677 30209 54711 30243
rect 54769 30209 54803 30243
rect 54953 30209 54987 30243
rect 55413 30209 55447 30243
rect 57161 30209 57195 30243
rect 57897 30209 57931 30243
rect 31125 30141 31159 30175
rect 38485 30141 38519 30175
rect 38761 30141 38795 30175
rect 42625 30141 42659 30175
rect 43637 30141 43671 30175
rect 50813 30141 50847 30175
rect 30665 30073 30699 30107
rect 39405 30073 39439 30107
rect 42809 30073 42843 30107
rect 1961 30005 1995 30039
rect 2513 30005 2547 30039
rect 26065 30005 26099 30039
rect 26433 30005 26467 30039
rect 29101 30005 29135 30039
rect 29469 30005 29503 30039
rect 31033 30005 31067 30039
rect 35265 30005 35299 30039
rect 36461 30005 36495 30039
rect 37657 30005 37691 30039
rect 38209 30005 38243 30039
rect 40325 30005 40359 30039
rect 40509 30005 40543 30039
rect 48145 30005 48179 30039
rect 57253 30005 57287 30039
rect 31125 29801 31159 29835
rect 38577 29801 38611 29835
rect 42441 29801 42475 29835
rect 43453 29801 43487 29835
rect 46949 29801 46983 29835
rect 47961 29801 47995 29835
rect 52101 29801 52135 29835
rect 54033 29801 54067 29835
rect 55413 29801 55447 29835
rect 31769 29733 31803 29767
rect 40233 29733 40267 29767
rect 27997 29665 28031 29699
rect 28089 29665 28123 29699
rect 31953 29665 31987 29699
rect 36737 29665 36771 29699
rect 39221 29665 39255 29699
rect 42165 29665 42199 29699
rect 45109 29665 45143 29699
rect 47685 29665 47719 29699
rect 51365 29665 51399 29699
rect 52745 29665 52779 29699
rect 53205 29665 53239 29699
rect 56517 29665 56551 29699
rect 57897 29665 57931 29699
rect 26893 29597 26927 29631
rect 27905 29597 27939 29631
rect 30849 29597 30883 29631
rect 31033 29597 31067 29631
rect 31677 29597 31711 29631
rect 33609 29597 33643 29631
rect 36093 29597 36127 29631
rect 37013 29597 37047 29631
rect 38761 29597 38795 29631
rect 38853 29597 38887 29631
rect 40049 29597 40083 29631
rect 40141 29597 40175 29631
rect 40325 29597 40359 29631
rect 40969 29597 41003 29631
rect 42073 29597 42107 29631
rect 43638 29591 43672 29625
rect 43821 29597 43855 29631
rect 44005 29597 44039 29631
rect 44097 29597 44131 29631
rect 45017 29597 45051 29631
rect 45201 29597 45235 29631
rect 46397 29597 46431 29631
rect 46765 29597 46799 29631
rect 47593 29597 47627 29631
rect 51273 29597 51307 29631
rect 51457 29597 51491 29631
rect 51917 29597 51951 29631
rect 52837 29597 52871 29631
rect 54217 29597 54251 29631
rect 54493 29597 54527 29631
rect 55321 29597 55355 29631
rect 55505 29597 55539 29631
rect 56333 29597 56367 29631
rect 27077 29529 27111 29563
rect 31217 29529 31251 29563
rect 33701 29529 33735 29563
rect 43729 29529 43763 29563
rect 46581 29529 46615 29563
rect 46673 29529 46707 29563
rect 27537 29461 27571 29495
rect 31953 29461 31987 29495
rect 36185 29461 36219 29495
rect 39037 29461 39071 29495
rect 39129 29461 39163 29495
rect 39865 29461 39899 29495
rect 41061 29461 41095 29495
rect 54401 29461 54435 29495
rect 28365 29257 28399 29291
rect 32505 29257 32539 29291
rect 42625 29257 42659 29291
rect 43361 29257 43395 29291
rect 43637 29257 43671 29291
rect 49985 29257 50019 29291
rect 50813 29257 50847 29291
rect 50997 29257 51031 29291
rect 51825 29257 51859 29291
rect 52745 29257 52779 29291
rect 54493 29257 54527 29291
rect 2145 29189 2179 29223
rect 33333 29189 33367 29223
rect 38577 29189 38611 29223
rect 40785 29189 40819 29223
rect 43269 29189 43303 29223
rect 1961 29121 1995 29155
rect 24593 29121 24627 29155
rect 26985 29121 27019 29155
rect 27252 29121 27286 29155
rect 30849 29121 30883 29155
rect 32137 29121 32171 29155
rect 37289 29121 37323 29155
rect 38485 29121 38519 29155
rect 38669 29121 38703 29155
rect 38853 29121 38887 29155
rect 38945 29121 38979 29155
rect 39405 29121 39439 29155
rect 40693 29121 40727 29155
rect 42533 29121 42567 29155
rect 42717 29121 42751 29155
rect 43177 29121 43211 29155
rect 43637 29121 43671 29155
rect 45937 29121 45971 29155
rect 46121 29121 46155 29155
rect 49893 29121 49927 29155
rect 50629 29121 50663 29155
rect 50905 29121 50939 29155
rect 51733 29121 51767 29155
rect 53113 29121 53147 29155
rect 54125 29121 54159 29155
rect 2789 29053 2823 29087
rect 24777 29053 24811 29087
rect 25329 29053 25363 29087
rect 31125 29053 31159 29087
rect 32229 29053 32263 29087
rect 37381 29053 37415 29087
rect 39681 29053 39715 29087
rect 43499 29053 43533 29087
rect 52929 29053 52963 29087
rect 53021 29053 53055 29087
rect 53205 29053 53239 29087
rect 54033 29053 54067 29087
rect 31033 28985 31067 29019
rect 33517 28985 33551 29019
rect 51181 28985 51215 29019
rect 30665 28917 30699 28951
rect 32321 28917 32355 28951
rect 37473 28917 37507 28951
rect 37657 28917 37691 28951
rect 38301 28917 38335 28951
rect 45937 28917 45971 28951
rect 25237 28713 25271 28747
rect 27169 28713 27203 28747
rect 48421 28713 48455 28747
rect 48789 28713 48823 28747
rect 52837 28713 52871 28747
rect 53573 28713 53607 28747
rect 54677 28713 54711 28747
rect 28825 28645 28859 28679
rect 29009 28645 29043 28679
rect 36921 28645 36955 28679
rect 41337 28645 41371 28679
rect 28549 28577 28583 28611
rect 29561 28577 29595 28611
rect 31309 28577 31343 28611
rect 34713 28577 34747 28611
rect 37565 28577 37599 28611
rect 51825 28577 51859 28611
rect 57805 28577 57839 28611
rect 25145 28509 25179 28543
rect 27169 28509 27203 28543
rect 27353 28509 27387 28543
rect 29837 28509 29871 28543
rect 31585 28509 31619 28543
rect 32689 28509 32723 28543
rect 32873 28509 32907 28543
rect 33425 28509 33459 28543
rect 33609 28509 33643 28543
rect 37749 28509 37783 28543
rect 38025 28509 38059 28543
rect 38853 28509 38887 28543
rect 39037 28509 39071 28543
rect 41153 28509 41187 28543
rect 43729 28509 43763 28543
rect 43913 28509 43947 28543
rect 45017 28509 45051 28543
rect 45165 28509 45199 28543
rect 45521 28509 45555 28543
rect 46673 28509 46707 28543
rect 46949 28509 46983 28543
rect 47593 28509 47627 28543
rect 47777 28509 47811 28543
rect 47869 28509 47903 28543
rect 48329 28509 48363 28543
rect 50169 28509 50203 28543
rect 50445 28509 50479 28543
rect 51457 28509 51491 28543
rect 52466 28509 52500 28543
rect 52929 28509 52963 28543
rect 54493 28509 54527 28543
rect 56333 28509 56367 28543
rect 32965 28441 32999 28475
rect 34980 28441 35014 28475
rect 36737 28441 36771 28475
rect 40325 28441 40359 28475
rect 40693 28441 40727 28475
rect 45293 28441 45327 28475
rect 45393 28441 45427 28475
rect 47409 28441 47443 28475
rect 51641 28441 51675 28475
rect 53481 28441 53515 28475
rect 54309 28441 54343 28475
rect 56517 28441 56551 28475
rect 33517 28373 33551 28407
rect 36093 28373 36127 28407
rect 37933 28373 37967 28407
rect 43913 28373 43947 28407
rect 45661 28373 45695 28407
rect 46489 28373 46523 28407
rect 46857 28373 46891 28407
rect 52285 28373 52319 28407
rect 52469 28373 52503 28407
rect 29015 28169 29049 28203
rect 33333 28169 33367 28203
rect 36461 28169 36495 28203
rect 43361 28169 43395 28203
rect 44373 28169 44407 28203
rect 44925 28169 44959 28203
rect 46029 28169 46063 28203
rect 47961 28169 47995 28203
rect 49617 28169 49651 28203
rect 50307 28169 50341 28203
rect 53941 28169 53975 28203
rect 54677 28169 54711 28203
rect 29101 28101 29135 28135
rect 30941 28101 30975 28135
rect 34060 28101 34094 28135
rect 41061 28101 41095 28135
rect 47593 28101 47627 28135
rect 51365 28101 51399 28135
rect 53230 28101 53264 28135
rect 47823 28067 47857 28101
rect 28917 28033 28951 28067
rect 29193 28033 29227 28067
rect 31217 28033 31251 28067
rect 31309 28033 31343 28067
rect 31401 28033 31435 28067
rect 31585 28033 31619 28067
rect 32137 28033 32171 28067
rect 33057 28033 33091 28067
rect 33793 28033 33827 28067
rect 35725 28033 35759 28067
rect 36369 28033 36403 28067
rect 36737 28033 36771 28067
rect 37289 28033 37323 28067
rect 37841 28033 37875 28067
rect 38025 28033 38059 28067
rect 38485 28033 38519 28067
rect 38577 28033 38611 28067
rect 39221 28033 39255 28067
rect 39405 28033 39439 28067
rect 43177 28033 43211 28067
rect 43361 28033 43395 28067
rect 44005 28033 44039 28067
rect 44833 28033 44867 28067
rect 45661 28033 45695 28067
rect 46489 28033 46523 28067
rect 46673 28033 46707 28067
rect 49433 28033 49467 28067
rect 49617 28033 49651 28067
rect 51549 28033 51583 28067
rect 51641 28033 51675 28067
rect 51917 28033 51951 28067
rect 52745 28033 52779 28067
rect 53849 28033 53883 28067
rect 54033 28033 54067 28067
rect 54493 28033 54527 28067
rect 54677 28033 54711 28067
rect 58081 28033 58115 28067
rect 29653 27965 29687 27999
rect 32229 27965 32263 27999
rect 33333 27965 33367 27999
rect 36553 27965 36587 27999
rect 39313 27965 39347 27999
rect 43913 27965 43947 27999
rect 45753 27965 45787 27999
rect 50077 27965 50111 27999
rect 53021 27965 53055 27999
rect 53113 27965 53147 27999
rect 29929 27897 29963 27931
rect 30113 27897 30147 27931
rect 33149 27897 33183 27931
rect 35817 27897 35851 27931
rect 51825 27897 51859 27931
rect 32137 27829 32171 27863
rect 32505 27829 32539 27863
rect 35173 27829 35207 27863
rect 36737 27829 36771 27863
rect 41153 27829 41187 27863
rect 46581 27829 46615 27863
rect 47777 27829 47811 27863
rect 53389 27829 53423 27863
rect 28825 27625 28859 27659
rect 32689 27625 32723 27659
rect 37105 27625 37139 27659
rect 37933 27625 37967 27659
rect 38117 27625 38151 27659
rect 38761 27625 38795 27659
rect 44005 27625 44039 27659
rect 46029 27625 46063 27659
rect 46397 27625 46431 27659
rect 47409 27625 47443 27659
rect 47961 27625 47995 27659
rect 52929 27625 52963 27659
rect 29009 27557 29043 27591
rect 33425 27557 33459 27591
rect 40693 27557 40727 27591
rect 45017 27557 45051 27591
rect 49617 27557 49651 27591
rect 56977 27557 57011 27591
rect 30941 27489 30975 27523
rect 31669 27489 31703 27523
rect 31861 27489 31895 27523
rect 31954 27489 31988 27523
rect 36277 27489 36311 27523
rect 36829 27489 36863 27523
rect 47501 27489 47535 27523
rect 50445 27489 50479 27523
rect 53573 27489 53607 27523
rect 2237 27421 2271 27455
rect 27997 27421 28031 27455
rect 28181 27421 28215 27455
rect 30481 27421 30515 27455
rect 30573 27421 30607 27455
rect 30849 27421 30883 27455
rect 31769 27421 31803 27455
rect 33333 27421 33367 27455
rect 33517 27421 33551 27455
rect 36185 27421 36219 27455
rect 36369 27421 36403 27455
rect 37105 27421 37139 27455
rect 37289 27421 37323 27455
rect 38577 27421 38611 27455
rect 41521 27421 41555 27455
rect 41797 27421 41831 27455
rect 42349 27421 42383 27455
rect 43637 27421 43671 27455
rect 45201 27421 45235 27455
rect 45477 27421 45511 27455
rect 45937 27421 45971 27455
rect 47225 27421 47259 27455
rect 47317 27421 47351 27455
rect 48145 27421 48179 27455
rect 48237 27421 48271 27455
rect 48421 27421 48455 27455
rect 48513 27421 48547 27455
rect 49065 27421 49099 27455
rect 49341 27421 49375 27455
rect 49433 27421 49467 27455
rect 50169 27421 50203 27455
rect 51457 27421 51491 27455
rect 51733 27421 51767 27455
rect 52745 27421 52779 27455
rect 53481 27421 53515 27455
rect 53665 27421 53699 27455
rect 56885 27421 56919 27455
rect 28641 27353 28675 27387
rect 28857 27353 28891 27387
rect 29837 27353 29871 27387
rect 32505 27353 32539 27387
rect 37749 27353 37783 27387
rect 37965 27353 37999 27387
rect 40509 27353 40543 27387
rect 41705 27353 41739 27387
rect 42533 27353 42567 27387
rect 43821 27353 43855 27387
rect 49249 27353 49283 27387
rect 28181 27285 28215 27319
rect 31493 27285 31527 27319
rect 32705 27285 32739 27319
rect 32873 27285 32907 27319
rect 41337 27285 41371 27319
rect 45385 27285 45419 27319
rect 32597 27081 32631 27115
rect 37749 27081 37783 27115
rect 46397 27081 46431 27115
rect 49249 27081 49283 27115
rect 51549 27081 51583 27115
rect 51825 27081 51859 27115
rect 57069 27081 57103 27115
rect 28733 27013 28767 27047
rect 32137 27013 32171 27047
rect 39497 27013 39531 27047
rect 41245 27013 41279 27047
rect 48881 27013 48915 27047
rect 49065 27013 49099 27047
rect 51089 27013 51123 27047
rect 1961 26945 1995 26979
rect 8769 26945 8803 26979
rect 28641 26945 28675 26979
rect 28825 26945 28859 26979
rect 29285 26945 29319 26979
rect 29469 26945 29503 26979
rect 31401 26945 31435 26979
rect 36553 26945 36587 26979
rect 36737 26945 36771 26979
rect 37565 26945 37599 26979
rect 37841 26945 37875 26979
rect 40141 26945 40175 26979
rect 40325 26945 40359 26979
rect 40877 26945 40911 26979
rect 41153 26945 41187 26979
rect 41429 26945 41463 26979
rect 43729 26945 43763 26979
rect 43913 26945 43947 26979
rect 46305 26945 46339 26979
rect 46765 26945 46799 26979
rect 48053 26945 48087 26979
rect 56885 26945 56919 26979
rect 2145 26877 2179 26911
rect 2789 26877 2823 26911
rect 9045 26877 9079 26911
rect 29929 26877 29963 26911
rect 30205 26877 30239 26911
rect 31217 26877 31251 26911
rect 36645 26877 36679 26911
rect 41705 26877 41739 26911
rect 49709 26877 49743 26911
rect 49985 26877 50019 26911
rect 51641 26877 51675 26911
rect 31585 26809 31619 26843
rect 32413 26809 32447 26843
rect 39681 26809 39715 26843
rect 51089 26809 51123 26843
rect 29285 26741 29319 26775
rect 37381 26741 37415 26775
rect 40141 26741 40175 26775
rect 43729 26741 43763 26775
rect 48145 26741 48179 26775
rect 58081 26741 58115 26775
rect 2513 26537 2547 26571
rect 47317 26537 47351 26571
rect 51273 26537 51307 26571
rect 51457 26537 51491 26571
rect 31585 26469 31619 26503
rect 40877 26469 40911 26503
rect 43269 26469 43303 26503
rect 43821 26469 43855 26503
rect 29837 26401 29871 26435
rect 30665 26401 30699 26435
rect 50445 26401 50479 26435
rect 56333 26401 56367 26435
rect 58173 26401 58207 26435
rect 2421 26333 2455 26367
rect 8953 26333 8987 26367
rect 9781 26333 9815 26367
rect 29745 26333 29779 26367
rect 29929 26333 29963 26367
rect 30389 26323 30423 26357
rect 30573 26333 30607 26367
rect 30757 26333 30791 26367
rect 30941 26333 30975 26367
rect 31769 26333 31803 26367
rect 31861 26333 31895 26367
rect 32045 26333 32079 26367
rect 32137 26333 32171 26367
rect 37565 26333 37599 26367
rect 37841 26333 37875 26367
rect 40049 26333 40083 26367
rect 40325 26333 40359 26367
rect 40785 26333 40819 26367
rect 41429 26333 41463 26367
rect 41613 26333 41647 26367
rect 43085 26333 43119 26367
rect 44005 26333 44039 26367
rect 44281 26333 44315 26367
rect 44465 26333 44499 26367
rect 47869 26333 47903 26367
rect 50169 26333 50203 26367
rect 50353 26333 50387 26367
rect 50573 26333 50607 26367
rect 37381 26265 37415 26299
rect 40233 26265 40267 26299
rect 41521 26265 41555 26299
rect 47225 26265 47259 26299
rect 50445 26265 50479 26299
rect 51089 26265 51123 26299
rect 51305 26265 51339 26299
rect 56517 26265 56551 26299
rect 31125 26197 31159 26231
rect 37749 26197 37783 26231
rect 39865 26197 39899 26231
rect 47961 26197 47995 26231
rect 41429 25993 41463 26027
rect 44741 25993 44775 26027
rect 57069 25993 57103 26027
rect 7757 25925 7791 25959
rect 8125 25857 8159 25891
rect 8769 25857 8803 25891
rect 30389 25857 30423 25891
rect 30481 25857 30515 25891
rect 30665 25857 30699 25891
rect 30757 25857 30791 25891
rect 31217 25857 31251 25891
rect 31401 25857 31435 25891
rect 37289 25857 37323 25891
rect 37565 25857 37599 25891
rect 37749 25857 37783 25891
rect 38025 25857 38059 25891
rect 38945 25857 38979 25891
rect 39773 25879 39807 25913
rect 39865 25891 39899 25925
rect 40003 25857 40037 25891
rect 40141 25857 40175 25891
rect 40233 25857 40267 25891
rect 40785 25857 40819 25891
rect 41613 25857 41647 25891
rect 41797 25857 41831 25891
rect 41889 25857 41923 25891
rect 43453 25857 43487 25891
rect 43637 25857 43671 25891
rect 43821 25857 43855 25891
rect 44465 25857 44499 25891
rect 48881 25857 48915 25891
rect 49065 25857 49099 25891
rect 56333 25857 56367 25891
rect 56977 25857 57011 25891
rect 9597 25789 9631 25823
rect 38761 25789 38795 25823
rect 38853 25789 38887 25823
rect 39037 25789 39071 25823
rect 44281 25789 44315 25823
rect 44833 25789 44867 25823
rect 37841 25721 37875 25755
rect 39589 25721 39623 25755
rect 30205 25653 30239 25687
rect 31217 25653 31251 25687
rect 38577 25653 38611 25687
rect 40877 25653 40911 25687
rect 49249 25653 49283 25687
rect 56425 25653 56459 25687
rect 58081 25653 58115 25687
rect 39313 25449 39347 25483
rect 44281 25449 44315 25483
rect 36829 25381 36863 25415
rect 40969 25381 41003 25415
rect 44465 25381 44499 25415
rect 36553 25313 36587 25347
rect 37381 25313 37415 25347
rect 40049 25313 40083 25347
rect 40224 25313 40258 25347
rect 56333 25313 56367 25347
rect 56517 25313 56551 25347
rect 58173 25313 58207 25347
rect 8953 25245 8987 25279
rect 36461 25245 36495 25279
rect 37473 25245 37507 25279
rect 38301 25245 38335 25279
rect 38485 25245 38519 25279
rect 38945 25245 38979 25279
rect 39129 25245 39163 25279
rect 40141 25245 40175 25279
rect 40325 25245 40359 25279
rect 41153 25245 41187 25279
rect 41797 25245 41831 25279
rect 42717 25245 42751 25279
rect 42809 25245 42843 25279
rect 42901 25245 42935 25279
rect 43085 25245 43119 25279
rect 45017 25245 45051 25279
rect 47133 25245 47167 25279
rect 47317 25245 47351 25279
rect 47777 25245 47811 25279
rect 47961 25245 47995 25279
rect 9873 25177 9907 25211
rect 40877 25177 40911 25211
rect 41061 25177 41095 25211
rect 41981 25177 42015 25211
rect 44097 25177 44131 25211
rect 37841 25109 37875 25143
rect 38485 25109 38519 25143
rect 39865 25109 39899 25143
rect 42441 25109 42475 25143
rect 44297 25109 44331 25143
rect 45201 25109 45235 25143
rect 47317 25109 47351 25143
rect 47869 25109 47903 25143
rect 38669 24905 38703 24939
rect 39431 24905 39465 24939
rect 44465 24905 44499 24939
rect 47961 24905 47995 24939
rect 37381 24837 37415 24871
rect 39221 24837 39255 24871
rect 41245 24837 41279 24871
rect 2329 24769 2363 24803
rect 8769 24769 8803 24803
rect 37565 24769 37599 24803
rect 37657 24769 37691 24803
rect 38485 24769 38519 24803
rect 38761 24769 38795 24803
rect 40233 24769 40267 24803
rect 41061 24769 41095 24803
rect 41337 24769 41371 24803
rect 41429 24769 41463 24803
rect 42625 24769 42659 24803
rect 42901 24769 42935 24803
rect 43453 24769 43487 24803
rect 45293 24769 45327 24803
rect 46508 24769 46542 24803
rect 46673 24769 46707 24803
rect 46765 24769 46799 24803
rect 47593 24769 47627 24803
rect 56885 24769 56919 24803
rect 9045 24701 9079 24735
rect 40325 24701 40359 24735
rect 44557 24701 44591 24735
rect 44649 24701 44683 24735
rect 47869 24701 47903 24735
rect 47961 24701 47995 24735
rect 37657 24633 37691 24667
rect 41613 24633 41647 24667
rect 42809 24633 42843 24667
rect 43637 24633 43671 24667
rect 46305 24633 46339 24667
rect 1869 24565 1903 24599
rect 2421 24565 2455 24599
rect 38485 24565 38519 24599
rect 39405 24565 39439 24599
rect 39589 24565 39623 24599
rect 40509 24565 40543 24599
rect 42441 24565 42475 24599
rect 44097 24565 44131 24599
rect 45385 24565 45419 24599
rect 45753 24565 45787 24599
rect 47685 24565 47719 24599
rect 56977 24565 57011 24599
rect 58081 24565 58115 24599
rect 40325 24361 40359 24395
rect 44465 24361 44499 24395
rect 46673 24361 46707 24395
rect 46213 24293 46247 24327
rect 32321 24225 32355 24259
rect 41429 24225 41463 24259
rect 44005 24225 44039 24259
rect 47225 24225 47259 24259
rect 47961 24225 47995 24259
rect 56333 24225 56367 24259
rect 56517 24225 56551 24259
rect 58173 24225 58207 24259
rect 39957 24157 39991 24191
rect 40141 24157 40175 24191
rect 41613 24157 41647 24191
rect 41889 24157 41923 24191
rect 42717 24157 42751 24191
rect 42809 24157 42843 24191
rect 42993 24157 43027 24191
rect 44097 24157 44131 24191
rect 45937 24157 45971 24191
rect 46029 24157 46063 24191
rect 48053 24157 48087 24191
rect 48881 24157 48915 24191
rect 32505 24089 32539 24123
rect 34161 24089 34195 24123
rect 41797 24089 41831 24123
rect 47041 24089 47075 24123
rect 49157 24089 49191 24123
rect 47133 24021 47167 24055
rect 48421 24021 48455 24055
rect 32597 23817 32631 23851
rect 43637 23817 43671 23851
rect 44097 23817 44131 23851
rect 45201 23817 45235 23851
rect 47961 23817 47995 23851
rect 2145 23749 2179 23783
rect 43545 23749 43579 23783
rect 44465 23749 44499 23783
rect 1961 23681 1995 23715
rect 32505 23681 32539 23715
rect 43361 23681 43395 23715
rect 43637 23681 43671 23715
rect 44281 23681 44315 23715
rect 44373 23681 44407 23715
rect 44649 23681 44683 23715
rect 44741 23681 44775 23715
rect 45477 23681 45511 23715
rect 45569 23681 45603 23715
rect 46673 23681 46707 23715
rect 46765 23681 46799 23715
rect 46857 23681 46891 23715
rect 47593 23681 47627 23715
rect 47777 23681 47811 23715
rect 2789 23613 2823 23647
rect 45385 23613 45419 23647
rect 45661 23613 45695 23647
rect 46581 23613 46615 23647
rect 46397 23545 46431 23579
rect 45017 23273 45051 23307
rect 47041 23273 47075 23307
rect 40417 23205 40451 23239
rect 40141 23137 40175 23171
rect 40969 23137 41003 23171
rect 41889 23137 41923 23171
rect 44097 23137 44131 23171
rect 45661 23137 45695 23171
rect 40049 23069 40083 23103
rect 41061 23069 41095 23103
rect 42073 23069 42107 23103
rect 42349 23069 42383 23103
rect 42993 23069 43027 23103
rect 43085 23069 43119 23103
rect 44281 23069 44315 23103
rect 46949 23069 46983 23103
rect 47133 23069 47167 23103
rect 42809 23001 42843 23035
rect 45385 23001 45419 23035
rect 41429 22933 41463 22967
rect 42257 22933 42291 22967
rect 43085 22933 43119 22967
rect 44465 22933 44499 22967
rect 45477 22933 45511 22967
rect 43729 22729 43763 22763
rect 44741 22729 44775 22763
rect 43361 22593 43395 22627
rect 43545 22593 43579 22627
rect 44373 22593 44407 22627
rect 45201 22593 45235 22627
rect 45385 22593 45419 22627
rect 56517 22593 56551 22627
rect 57161 22593 57195 22627
rect 44465 22525 44499 22559
rect 45293 22525 45327 22559
rect 56609 22389 56643 22423
rect 57253 22389 57287 22423
rect 58081 22389 58115 22423
rect 43545 22185 43579 22219
rect 44189 22185 44223 22219
rect 56333 22049 56367 22083
rect 56517 22049 56551 22083
rect 57897 22049 57931 22083
rect 2237 21981 2271 22015
rect 44465 21981 44499 22015
rect 43361 21913 43395 21947
rect 43566 21913 43600 21947
rect 44189 21913 44223 21947
rect 43729 21845 43763 21879
rect 44373 21845 44407 21879
rect 17141 21641 17175 21675
rect 1961 21505 1995 21539
rect 17049 21505 17083 21539
rect 19625 21505 19659 21539
rect 29745 21505 29779 21539
rect 56977 21505 57011 21539
rect 2145 21437 2179 21471
rect 2789 21437 2823 21471
rect 20177 21437 20211 21471
rect 31493 21437 31527 21471
rect 57069 21301 57103 21335
rect 58081 21301 58115 21335
rect 31309 20961 31343 20995
rect 56333 20961 56367 20995
rect 57897 20961 57931 20995
rect 2237 20893 2271 20927
rect 18429 20893 18463 20927
rect 19625 20893 19659 20927
rect 28641 20893 28675 20927
rect 30481 20893 30515 20927
rect 20177 20825 20211 20859
rect 29009 20825 29043 20859
rect 56517 20825 56551 20859
rect 18613 20757 18647 20791
rect 30573 20485 30607 20519
rect 1961 20417 1995 20451
rect 19533 20417 19567 20451
rect 29653 20417 29687 20451
rect 58081 20417 58115 20451
rect 2145 20349 2179 20383
rect 2789 20349 2823 20383
rect 20361 20349 20395 20383
rect 2605 20009 2639 20043
rect 31125 19873 31159 19907
rect 56333 19873 56367 19907
rect 56517 19873 56551 19907
rect 57805 19873 57839 19907
rect 2513 19805 2547 19839
rect 19533 19805 19567 19839
rect 30481 19805 30515 19839
rect 20453 19737 20487 19771
rect 2513 19465 2547 19499
rect 2421 19329 2455 19363
rect 19533 19329 19567 19363
rect 20085 19329 20119 19363
rect 29561 19329 29595 19363
rect 29837 19329 29871 19363
rect 2513 18717 2547 18751
rect 3801 18717 3835 18751
rect 3893 18581 3927 18615
rect 2421 18309 2455 18343
rect 2237 18241 2271 18275
rect 30389 18241 30423 18275
rect 2789 18173 2823 18207
rect 30481 18037 30515 18071
rect 58081 18037 58115 18071
rect 31033 17697 31067 17731
rect 31217 17697 31251 17731
rect 56333 17697 56367 17731
rect 58173 17697 58207 17731
rect 2237 17629 2271 17663
rect 32873 17561 32907 17595
rect 56517 17561 56551 17595
rect 57161 17289 57195 17323
rect 1961 17153 1995 17187
rect 57069 17153 57103 17187
rect 2145 17085 2179 17119
rect 2789 17085 2823 17119
rect 58081 16949 58115 16983
rect 2421 16745 2455 16779
rect 56333 16609 56367 16643
rect 57805 16609 57839 16643
rect 2329 16541 2363 16575
rect 56517 16473 56551 16507
rect 57161 16201 57195 16235
rect 57069 16065 57103 16099
rect 58081 15861 58115 15895
rect 56333 15521 56367 15555
rect 57897 15521 57931 15555
rect 56517 15385 56551 15419
rect 56977 15113 57011 15147
rect 56885 14977 56919 15011
rect 58081 14773 58115 14807
rect 56333 14433 56367 14467
rect 2237 14365 2271 14399
rect 56517 14297 56551 14331
rect 58173 14297 58207 14331
rect 56977 14025 57011 14059
rect 1961 13889 1995 13923
rect 56885 13889 56919 13923
rect 2145 13821 2179 13855
rect 2789 13821 2823 13855
rect 2513 13481 2547 13515
rect 2421 13277 2455 13311
rect 1777 12733 1811 12767
rect 2237 12733 2271 12767
rect 2421 12733 2455 12767
rect 3985 12733 4019 12767
rect 3893 12393 3927 12427
rect 2237 12189 2271 12223
rect 3801 12189 3835 12223
rect 1961 11713 1995 11747
rect 2145 11645 2179 11679
rect 2789 11645 2823 11679
rect 2421 11305 2455 11339
rect 2329 11101 2363 11135
rect 30021 10081 30055 10115
rect 57989 10081 58023 10115
rect 29561 10013 29595 10047
rect 56609 10013 56643 10047
rect 29745 9945 29779 9979
rect 57253 9945 57287 9979
rect 56701 9877 56735 9911
rect 29653 9673 29687 9707
rect 29561 9537 29595 9571
rect 58081 9333 58115 9367
rect 56333 8993 56367 9027
rect 56517 8993 56551 9027
rect 57897 8993 57931 9027
rect 2237 8925 2271 8959
rect 1961 8449 1995 8483
rect 2145 8381 2179 8415
rect 2789 8381 2823 8415
rect 2145 8041 2179 8075
rect 1593 7837 1627 7871
rect 2053 7837 2087 7871
rect 2697 7837 2731 7871
rect 2789 7701 2823 7735
rect 2145 7429 2179 7463
rect 1961 7361 1995 7395
rect 4261 7361 4295 7395
rect 2789 7293 2823 7327
rect 4353 7157 4387 7191
rect 1409 6817 1443 6851
rect 3985 6817 4019 6851
rect 56977 6749 57011 6783
rect 57805 6749 57839 6783
rect 1593 6681 1627 6715
rect 3249 6681 3283 6715
rect 57069 6613 57103 6647
rect 5181 6341 5215 6375
rect 4261 6273 4295 6307
rect 55597 6273 55631 6307
rect 57897 6273 57931 6307
rect 1961 6205 1995 6239
rect 2145 6205 2179 6239
rect 2881 6205 2915 6239
rect 56885 6069 56919 6103
rect 57989 6069 58023 6103
rect 1869 5865 1903 5899
rect 2421 5865 2455 5899
rect 56333 5729 56367 5763
rect 56517 5729 56551 5763
rect 58173 5729 58207 5763
rect 2329 5661 2363 5695
rect 2973 5661 3007 5695
rect 55873 5661 55907 5695
rect 3065 5525 3099 5559
rect 2145 5253 2179 5287
rect 55689 5253 55723 5287
rect 55505 5185 55539 5219
rect 1961 5117 1995 5151
rect 2789 5117 2823 5151
rect 57345 5117 57379 5151
rect 8309 4981 8343 5015
rect 58081 4981 58115 5015
rect 1869 4777 1903 4811
rect 56333 4641 56367 4675
rect 56793 4641 56827 4675
rect 2513 4573 2547 4607
rect 7849 4573 7883 4607
rect 9137 4573 9171 4607
rect 54769 4573 54803 4607
rect 55873 4573 55907 4607
rect 56517 4505 56551 4539
rect 7941 4437 7975 4471
rect 9229 4437 9263 4471
rect 8217 4165 8251 4199
rect 2237 4097 2271 4131
rect 7389 4097 7423 4131
rect 14841 4097 14875 4131
rect 22477 4097 22511 4131
rect 26985 4097 27019 4131
rect 31125 4097 31159 4131
rect 38025 4097 38059 4131
rect 49985 4097 50019 4131
rect 53849 4097 53883 4131
rect 54861 4097 54895 4131
rect 55505 4097 55539 4131
rect 57897 4097 57931 4131
rect 2421 4029 2455 4063
rect 2789 4029 2823 4063
rect 8033 4029 8067 4063
rect 8493 4029 8527 4063
rect 55703 4029 55737 4063
rect 57345 4029 57379 4063
rect 57989 3961 58023 3995
rect 4721 3893 4755 3927
rect 7481 3893 7515 3927
rect 14933 3893 14967 3927
rect 16865 3893 16899 3927
rect 22569 3893 22603 3927
rect 23305 3893 23339 3927
rect 27077 3893 27111 3927
rect 30021 3893 30055 3927
rect 30665 3893 30699 3927
rect 31217 3893 31251 3927
rect 32321 3893 32355 3927
rect 38117 3893 38151 3927
rect 46489 3893 46523 3927
rect 50077 3893 50111 3927
rect 53941 3893 53975 3927
rect 54953 3893 54987 3927
rect 1869 3689 1903 3723
rect 3801 3553 3835 3587
rect 4261 3553 4295 3587
rect 6561 3553 6595 3587
rect 9597 3553 9631 3587
rect 9873 3553 9907 3587
rect 15301 3553 15335 3587
rect 20821 3553 20855 3587
rect 25145 3553 25179 3587
rect 26893 3553 26927 3587
rect 27169 3553 27203 3587
rect 29837 3553 29871 3587
rect 32137 3553 32171 3587
rect 32873 3553 32907 3587
rect 46305 3553 46339 3587
rect 47041 3553 47075 3587
rect 50353 3553 50387 3587
rect 50629 3553 50663 3587
rect 53113 3553 53147 3587
rect 54125 3553 54159 3587
rect 56333 3553 56367 3587
rect 57897 3553 57931 3587
rect 1777 3485 1811 3519
rect 2421 3485 2455 3519
rect 3065 3485 3099 3519
rect 6101 3485 6135 3519
rect 9413 3485 9447 3519
rect 12265 3485 12299 3519
rect 13093 3485 13127 3519
rect 15117 3485 15151 3519
rect 17417 3485 17451 3519
rect 19717 3485 19751 3519
rect 20361 3485 20395 3519
rect 22845 3485 22879 3519
rect 23857 3485 23891 3519
rect 24409 3485 24443 3519
rect 26709 3485 26743 3519
rect 38577 3485 38611 3519
rect 48789 3485 48823 3519
rect 49617 3485 49651 3519
rect 50169 3485 50203 3519
rect 52929 3485 52963 3519
rect 55321 3485 55355 3519
rect 3157 3417 3191 3451
rect 3985 3417 4019 3451
rect 6285 3417 6319 3451
rect 16957 3417 16991 3451
rect 19809 3417 19843 3451
rect 20545 3417 20579 3451
rect 22937 3417 22971 3451
rect 24593 3417 24627 3451
rect 30021 3417 30055 3451
rect 31677 3417 31711 3451
rect 32321 3417 32355 3451
rect 46489 3417 46523 3451
rect 56517 3417 56551 3451
rect 2513 3349 2547 3383
rect 12357 3349 12391 3383
rect 17509 3349 17543 3383
rect 55413 3349 55447 3383
rect 4629 3145 4663 3179
rect 32689 3145 32723 3179
rect 46857 3145 46891 3179
rect 56977 3145 57011 3179
rect 57989 3145 58023 3179
rect 2329 3077 2363 3111
rect 12725 3077 12759 3111
rect 16865 3077 16899 3111
rect 23029 3077 23063 3111
rect 29929 3077 29963 3111
rect 38485 3077 38519 3111
rect 47685 3077 47719 3111
rect 48421 3077 48455 3111
rect 54217 3077 54251 3111
rect 4537 3009 4571 3043
rect 5365 3009 5399 3043
rect 12541 3009 12575 3043
rect 15393 3009 15427 3043
rect 16681 3009 16715 3043
rect 20545 3009 20579 3043
rect 22845 3009 22879 3043
rect 27169 3009 27203 3043
rect 29745 3009 29779 3043
rect 32597 3009 32631 3043
rect 38301 3009 38335 3043
rect 46765 3009 46799 3043
rect 47593 3009 47627 3043
rect 48237 3009 48271 3043
rect 53573 3009 53607 3043
rect 56885 3009 56919 3043
rect 57897 3009 57931 3043
rect 2145 2941 2179 2975
rect 2605 2941 2639 2975
rect 7573 2941 7607 2975
rect 8033 2941 8067 2975
rect 8217 2941 8251 2975
rect 9137 2941 9171 2975
rect 13001 2941 13035 2975
rect 17141 2941 17175 2975
rect 23305 2941 23339 2975
rect 30941 2941 30975 2975
rect 38761 2941 38795 2975
rect 49617 2941 49651 2975
rect 54033 2941 54067 2975
rect 54769 2941 54803 2975
rect 6929 2805 6963 2839
rect 2421 2601 2455 2635
rect 9045 2601 9079 2635
rect 9781 2601 9815 2635
rect 31217 2601 31251 2635
rect 54217 2601 54251 2635
rect 58081 2601 58115 2635
rect 6561 2465 6595 2499
rect 7021 2465 7055 2499
rect 55505 2465 55539 2499
rect 8953 2397 8987 2431
rect 31125 2397 31159 2431
rect 6745 2329 6779 2363
rect 55689 2329 55723 2363
rect 57345 2329 57379 2363
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 658 57400 664 57452
rect 716 57440 722 57452
rect 1397 57443 1455 57449
rect 1397 57440 1409 57443
rect 716 57412 1409 57440
rect 716 57400 722 57412
rect 1397 57409 1409 57412
rect 1443 57409 1455 57443
rect 1397 57403 1455 57409
rect 10318 57400 10324 57452
rect 10376 57440 10382 57452
rect 10597 57443 10655 57449
rect 10597 57440 10609 57443
rect 10376 57412 10609 57440
rect 10376 57400 10382 57412
rect 10597 57409 10609 57412
rect 10643 57409 10655 57443
rect 10597 57403 10655 57409
rect 33502 57400 33508 57452
rect 33560 57440 33566 57452
rect 33781 57443 33839 57449
rect 33781 57440 33793 57443
rect 33560 57412 33793 57440
rect 33560 57400 33566 57412
rect 33781 57409 33793 57412
rect 33827 57409 33839 57443
rect 33781 57403 33839 57409
rect 57149 57443 57207 57449
rect 57149 57409 57161 57443
rect 57195 57440 57207 57443
rect 57698 57440 57704 57452
rect 57195 57412 57704 57440
rect 57195 57409 57207 57412
rect 57149 57403 57207 57409
rect 57698 57400 57704 57412
rect 57756 57400 57762 57452
rect 1673 57375 1731 57381
rect 1673 57341 1685 57375
rect 1719 57372 1731 57375
rect 20438 57372 20444 57384
rect 1719 57344 20444 57372
rect 1719 57341 1731 57344
rect 1673 57335 1731 57341
rect 20438 57332 20444 57344
rect 20496 57332 20502 57384
rect 10413 57307 10471 57313
rect 10413 57273 10425 57307
rect 10459 57304 10471 57307
rect 22002 57304 22008 57316
rect 10459 57276 22008 57304
rect 10459 57273 10471 57276
rect 10413 57267 10471 57273
rect 22002 57264 22008 57276
rect 22060 57264 22066 57316
rect 2869 57239 2927 57245
rect 2869 57205 2881 57239
rect 2915 57236 2927 57239
rect 3694 57236 3700 57248
rect 2915 57208 3700 57236
rect 2915 57205 2927 57208
rect 2869 57199 2927 57205
rect 3694 57196 3700 57208
rect 3752 57196 3758 57248
rect 3786 57196 3792 57248
rect 3844 57236 3850 57248
rect 4065 57239 4123 57245
rect 4065 57236 4077 57239
rect 3844 57208 4077 57236
rect 3844 57196 3850 57208
rect 4065 57205 4077 57208
rect 4111 57205 4123 57239
rect 17954 57236 17960 57248
rect 17915 57208 17960 57236
rect 4065 57199 4123 57205
rect 17954 57196 17960 57208
rect 18012 57196 18018 57248
rect 18046 57196 18052 57248
rect 18104 57236 18110 57248
rect 19242 57236 19248 57248
rect 18104 57208 19248 57236
rect 18104 57196 18110 57208
rect 19242 57196 19248 57208
rect 19300 57196 19306 57248
rect 31294 57196 31300 57248
rect 31352 57236 31358 57248
rect 31481 57239 31539 57245
rect 31481 57236 31493 57239
rect 31352 57208 31493 57236
rect 31352 57196 31358 57208
rect 31481 57205 31493 57208
rect 31527 57205 31539 57239
rect 31481 57199 31539 57205
rect 32122 57196 32128 57248
rect 32180 57236 32186 57248
rect 32309 57239 32367 57245
rect 32309 57236 32321 57239
rect 32180 57208 32321 57236
rect 32180 57196 32186 57208
rect 32309 57205 32321 57208
rect 32355 57205 32367 57239
rect 33594 57236 33600 57248
rect 33555 57208 33600 57236
rect 32309 57199 32367 57205
rect 33594 57196 33600 57208
rect 33652 57196 33658 57248
rect 35618 57196 35624 57248
rect 35676 57236 35682 57248
rect 35897 57239 35955 57245
rect 35897 57236 35909 57239
rect 35676 57208 35909 57236
rect 35676 57196 35682 57208
rect 35897 57205 35909 57208
rect 35943 57205 35955 57239
rect 35897 57199 35955 57205
rect 56045 57239 56103 57245
rect 56045 57205 56057 57239
rect 56091 57236 56103 57239
rect 56318 57236 56324 57248
rect 56091 57208 56324 57236
rect 56091 57205 56103 57208
rect 56045 57199 56103 57205
rect 56318 57196 56324 57208
rect 56376 57196 56382 57248
rect 56594 57196 56600 57248
rect 56652 57236 56658 57248
rect 56689 57239 56747 57245
rect 56689 57236 56701 57239
rect 56652 57208 56701 57236
rect 56652 57196 56658 57208
rect 56689 57205 56701 57208
rect 56735 57205 56747 57239
rect 57238 57236 57244 57248
rect 57199 57208 57244 57236
rect 56689 57199 56747 57205
rect 57238 57196 57244 57208
rect 57296 57196 57302 57248
rect 57422 57196 57428 57248
rect 57480 57236 57486 57248
rect 58069 57239 58127 57245
rect 58069 57236 58081 57239
rect 57480 57208 58081 57236
rect 57480 57196 57486 57208
rect 58069 57205 58081 57208
rect 58115 57205 58127 57239
rect 58069 57199 58127 57205
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 3786 56896 3792 56908
rect 3747 56868 3792 56896
rect 3786 56856 3792 56868
rect 3844 56856 3850 56908
rect 4154 56856 4160 56908
rect 4212 56896 4218 56908
rect 4249 56899 4307 56905
rect 4249 56896 4261 56899
rect 4212 56868 4261 56896
rect 4212 56856 4218 56868
rect 4249 56865 4261 56868
rect 4295 56865 4307 56899
rect 46658 56896 46664 56908
rect 4249 56859 4307 56865
rect 17420 56868 46664 56896
rect 1946 56788 1952 56840
rect 2004 56828 2010 56840
rect 2225 56831 2283 56837
rect 2225 56828 2237 56831
rect 2004 56800 2237 56828
rect 2004 56788 2010 56800
rect 2225 56797 2237 56800
rect 2271 56797 2283 56831
rect 2866 56828 2872 56840
rect 2827 56800 2872 56828
rect 2225 56791 2283 56797
rect 2866 56788 2872 56800
rect 2924 56788 2930 56840
rect 6362 56788 6368 56840
rect 6420 56828 6426 56840
rect 6457 56831 6515 56837
rect 6457 56828 6469 56831
rect 6420 56800 6469 56828
rect 6420 56788 6426 56800
rect 6457 56797 6469 56800
rect 6503 56797 6515 56831
rect 6457 56791 6515 56797
rect 7653 56831 7711 56837
rect 7653 56797 7665 56831
rect 7699 56828 7711 56831
rect 8662 56828 8668 56840
rect 7699 56800 8668 56828
rect 7699 56797 7711 56800
rect 7653 56791 7711 56797
rect 8662 56788 8668 56800
rect 8720 56788 8726 56840
rect 13262 56788 13268 56840
rect 13320 56828 13326 56840
rect 13449 56831 13507 56837
rect 13449 56828 13461 56831
rect 13320 56800 13461 56828
rect 13320 56788 13326 56800
rect 13449 56797 13461 56800
rect 13495 56797 13507 56831
rect 16022 56828 16028 56840
rect 15983 56800 16028 56828
rect 13449 56791 13507 56797
rect 16022 56788 16028 56800
rect 16080 56788 16086 56840
rect 17310 56788 17316 56840
rect 17368 56828 17374 56840
rect 17420 56837 17448 56868
rect 46658 56856 46664 56868
rect 46716 56856 46722 56908
rect 56318 56896 56324 56908
rect 56279 56868 56324 56896
rect 56318 56856 56324 56868
rect 56376 56856 56382 56908
rect 57974 56896 57980 56908
rect 57935 56868 57980 56896
rect 57974 56856 57980 56868
rect 58032 56856 58038 56908
rect 17405 56831 17463 56837
rect 17405 56828 17417 56831
rect 17368 56800 17417 56828
rect 17368 56788 17374 56800
rect 17405 56797 17417 56800
rect 17451 56797 17463 56831
rect 18230 56828 18236 56840
rect 18191 56800 18236 56828
rect 17405 56791 17463 56797
rect 18230 56788 18236 56800
rect 18288 56788 18294 56840
rect 22554 56828 22560 56840
rect 22515 56800 22560 56828
rect 22554 56788 22560 56800
rect 22612 56788 22618 56840
rect 27246 56828 27252 56840
rect 27207 56800 27252 56828
rect 27246 56788 27252 56800
rect 27304 56788 27310 56840
rect 27890 56828 27896 56840
rect 27851 56800 27896 56828
rect 27890 56788 27896 56800
rect 27948 56788 27954 56840
rect 28258 56788 28264 56840
rect 28316 56828 28322 56840
rect 28353 56831 28411 56837
rect 28353 56828 28365 56831
rect 28316 56800 28365 56828
rect 28316 56788 28322 56800
rect 28353 56797 28365 56800
rect 28399 56797 28411 56831
rect 30190 56828 30196 56840
rect 30151 56800 30196 56828
rect 28353 56791 28411 56797
rect 30190 56788 30196 56800
rect 30248 56788 30254 56840
rect 30650 56828 30656 56840
rect 30611 56800 30656 56828
rect 30650 56788 30656 56800
rect 30708 56788 30714 56840
rect 31294 56828 31300 56840
rect 31255 56800 31300 56828
rect 31294 56788 31300 56800
rect 31352 56788 31358 56840
rect 35618 56828 35624 56840
rect 35579 56800 35624 56828
rect 35618 56788 35624 56800
rect 35676 56788 35682 56840
rect 40034 56828 40040 56840
rect 39995 56800 40040 56828
rect 40034 56788 40040 56800
rect 40092 56788 40098 56840
rect 42242 56828 42248 56840
rect 42203 56800 42248 56828
rect 42242 56788 42248 56800
rect 42300 56788 42306 56840
rect 42886 56828 42892 56840
rect 42847 56800 42892 56828
rect 42886 56788 42892 56800
rect 42944 56788 42950 56840
rect 46198 56788 46204 56840
rect 46256 56828 46262 56840
rect 46477 56831 46535 56837
rect 46477 56828 46489 56831
rect 46256 56800 46489 56828
rect 46256 56788 46262 56800
rect 46477 56797 46489 56800
rect 46523 56797 46535 56831
rect 46477 56791 46535 56797
rect 49694 56788 49700 56840
rect 49752 56828 49758 56840
rect 50341 56831 50399 56837
rect 50341 56828 50353 56831
rect 49752 56800 50353 56828
rect 49752 56788 49758 56800
rect 50341 56797 50353 56800
rect 50387 56797 50399 56831
rect 50341 56791 50399 56797
rect 55490 56788 55496 56840
rect 55548 56828 55554 56840
rect 55861 56831 55919 56837
rect 55861 56828 55873 56831
rect 55548 56800 55873 56828
rect 55548 56788 55554 56800
rect 55861 56797 55873 56800
rect 55907 56797 55919 56831
rect 55861 56791 55919 56797
rect 3973 56763 4031 56769
rect 3973 56729 3985 56763
rect 4019 56760 4031 56763
rect 4338 56760 4344 56772
rect 4019 56732 4344 56760
rect 4019 56729 4031 56732
rect 3973 56723 4031 56729
rect 4338 56720 4344 56732
rect 4396 56720 4402 56772
rect 30745 56763 30803 56769
rect 30745 56729 30757 56763
rect 30791 56760 30803 56763
rect 31481 56763 31539 56769
rect 31481 56760 31493 56763
rect 30791 56732 31493 56760
rect 30791 56729 30803 56732
rect 30745 56723 30803 56729
rect 31481 56729 31493 56732
rect 31527 56729 31539 56763
rect 31481 56723 31539 56729
rect 31754 56720 31760 56772
rect 31812 56760 31818 56772
rect 33137 56763 33195 56769
rect 33137 56760 33149 56763
rect 31812 56732 33149 56760
rect 31812 56720 31818 56732
rect 33137 56729 33149 56732
rect 33183 56729 33195 56763
rect 35802 56760 35808 56772
rect 35763 56732 35808 56760
rect 33137 56723 33195 56729
rect 35802 56720 35808 56732
rect 35860 56720 35866 56772
rect 36078 56720 36084 56772
rect 36136 56760 36142 56772
rect 37461 56763 37519 56769
rect 37461 56760 37473 56763
rect 36136 56732 37473 56760
rect 36136 56720 36142 56732
rect 37461 56729 37473 56732
rect 37507 56729 37519 56763
rect 37461 56723 37519 56729
rect 56505 56763 56563 56769
rect 56505 56729 56517 56763
rect 56551 56760 56563 56763
rect 57974 56760 57980 56772
rect 56551 56732 57980 56760
rect 56551 56729 56563 56732
rect 56505 56723 56563 56729
rect 57974 56720 57980 56732
rect 58032 56720 58038 56772
rect 17497 56695 17555 56701
rect 17497 56661 17509 56695
rect 17543 56692 17555 56695
rect 17862 56692 17868 56704
rect 17543 56664 17868 56692
rect 17543 56661 17555 56664
rect 17497 56655 17555 56661
rect 17862 56652 17868 56664
rect 17920 56652 17926 56704
rect 22370 56692 22376 56704
rect 22331 56664 22376 56692
rect 22370 56652 22376 56664
rect 22428 56652 22434 56704
rect 27065 56695 27123 56701
rect 27065 56661 27077 56695
rect 27111 56692 27123 56695
rect 27154 56692 27160 56704
rect 27111 56664 27160 56692
rect 27111 56661 27123 56664
rect 27065 56655 27123 56661
rect 27154 56652 27160 56664
rect 27212 56652 27218 56704
rect 28166 56652 28172 56704
rect 28224 56692 28230 56704
rect 28445 56695 28503 56701
rect 28445 56692 28457 56695
rect 28224 56664 28457 56692
rect 28224 56652 28230 56664
rect 28445 56661 28457 56664
rect 28491 56661 28503 56695
rect 28445 56655 28503 56661
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 4338 56488 4344 56500
rect 4299 56460 4344 56488
rect 4338 56448 4344 56460
rect 4396 56448 4402 56500
rect 22189 56491 22247 56497
rect 22189 56457 22201 56491
rect 22235 56488 22247 56491
rect 22554 56488 22560 56500
rect 22235 56460 22560 56488
rect 22235 56457 22247 56460
rect 22189 56451 22247 56457
rect 22554 56448 22560 56460
rect 22612 56448 22618 56500
rect 24397 56491 24455 56497
rect 24397 56457 24409 56491
rect 24443 56488 24455 56491
rect 26970 56488 26976 56500
rect 24443 56460 26976 56488
rect 24443 56457 24455 56460
rect 24397 56451 24455 56457
rect 26970 56448 26976 56460
rect 27028 56448 27034 56500
rect 27246 56448 27252 56500
rect 27304 56488 27310 56500
rect 27341 56491 27399 56497
rect 27341 56488 27353 56491
rect 27304 56460 27353 56488
rect 27304 56448 27310 56460
rect 27341 56457 27353 56460
rect 27387 56457 27399 56491
rect 47854 56488 47860 56500
rect 27341 56451 27399 56457
rect 35866 56460 47860 56488
rect 18230 56420 18236 56432
rect 16776 56392 18236 56420
rect 1946 56352 1952 56364
rect 1907 56324 1952 56352
rect 1946 56312 1952 56324
rect 2004 56312 2010 56364
rect 4249 56355 4307 56361
rect 4249 56321 4261 56355
rect 4295 56321 4307 56355
rect 6362 56352 6368 56364
rect 6323 56324 6368 56352
rect 4249 56315 4307 56321
rect 2130 56284 2136 56296
rect 2091 56256 2136 56284
rect 2130 56244 2136 56256
rect 2188 56244 2194 56296
rect 2774 56284 2780 56296
rect 2735 56256 2780 56284
rect 2774 56244 2780 56256
rect 2832 56244 2838 56296
rect 4264 56148 4292 56315
rect 6362 56312 6368 56324
rect 6420 56312 6426 56364
rect 8662 56352 8668 56364
rect 8623 56324 8668 56352
rect 8662 56312 8668 56324
rect 8720 56312 8726 56364
rect 13262 56352 13268 56364
rect 13223 56324 13268 56352
rect 13262 56312 13268 56324
rect 13320 56312 13326 56364
rect 16776 56361 16804 56392
rect 18230 56380 18236 56392
rect 18288 56380 18294 56432
rect 22370 56380 22376 56432
rect 22428 56420 22434 56432
rect 23262 56423 23320 56429
rect 23262 56420 23274 56423
rect 22428 56392 23274 56420
rect 22428 56380 22434 56392
rect 23262 56389 23274 56392
rect 23308 56389 23320 56423
rect 28166 56420 28172 56432
rect 28127 56392 28172 56420
rect 23262 56383 23320 56389
rect 28166 56380 28172 56392
rect 28224 56380 28230 56432
rect 30650 56380 30656 56432
rect 30708 56420 30714 56432
rect 31478 56420 31484 56432
rect 30708 56392 31484 56420
rect 30708 56380 30714 56392
rect 16761 56355 16819 56361
rect 16761 56321 16773 56355
rect 16807 56321 16819 56355
rect 22002 56352 22008 56364
rect 21963 56324 22008 56352
rect 16761 56315 16819 56321
rect 22002 56312 22008 56324
rect 22060 56312 22066 56364
rect 26142 56312 26148 56364
rect 26200 56352 26206 56364
rect 26237 56355 26295 56361
rect 26237 56352 26249 56355
rect 26200 56324 26249 56352
rect 26200 56312 26206 56324
rect 26237 56321 26249 56324
rect 26283 56352 26295 56355
rect 27157 56355 27215 56361
rect 27157 56352 27169 56355
rect 26283 56324 27169 56352
rect 26283 56321 26295 56324
rect 26237 56315 26295 56321
rect 27157 56321 27169 56324
rect 27203 56321 27215 56355
rect 27157 56315 27215 56321
rect 27890 56312 27896 56364
rect 27948 56352 27954 56364
rect 30852 56361 30880 56392
rect 31478 56380 31484 56392
rect 31536 56420 31542 56432
rect 35866 56420 35894 56460
rect 47854 56448 47860 56460
rect 47912 56448 47918 56500
rect 40034 56420 40040 56432
rect 31536 56392 35894 56420
rect 39684 56392 40040 56420
rect 31536 56380 31542 56392
rect 27985 56355 28043 56361
rect 27985 56352 27997 56355
rect 27948 56324 27997 56352
rect 27948 56312 27954 56324
rect 27985 56321 27997 56324
rect 28031 56321 28043 56355
rect 27985 56315 28043 56321
rect 30837 56355 30895 56361
rect 30837 56321 30849 56355
rect 30883 56321 30895 56355
rect 32122 56352 32128 56364
rect 32083 56324 32128 56352
rect 30837 56315 30895 56321
rect 32122 56312 32128 56324
rect 32180 56312 32186 56364
rect 39684 56361 39712 56392
rect 40034 56380 40040 56392
rect 40092 56380 40098 56432
rect 42886 56420 42892 56432
rect 42628 56392 42892 56420
rect 42628 56361 42656 56392
rect 42886 56380 42892 56392
rect 42944 56380 42950 56432
rect 44450 56420 44456 56432
rect 44411 56392 44456 56420
rect 44450 56380 44456 56392
rect 44508 56380 44514 56432
rect 49694 56420 49700 56432
rect 49528 56392 49700 56420
rect 39669 56355 39727 56361
rect 39669 56321 39681 56355
rect 39715 56321 39727 56355
rect 39669 56315 39727 56321
rect 42613 56355 42671 56361
rect 42613 56321 42625 56355
rect 42659 56321 42671 56355
rect 46658 56352 46664 56364
rect 46619 56324 46664 56352
rect 42613 56315 42671 56321
rect 46658 56312 46664 56324
rect 46716 56312 46722 56364
rect 49528 56361 49556 56392
rect 49694 56380 49700 56392
rect 49752 56380 49758 56432
rect 55677 56423 55735 56429
rect 55677 56389 55689 56423
rect 55723 56420 55735 56423
rect 57977 56423 58035 56429
rect 57977 56420 57989 56423
rect 55723 56392 57989 56420
rect 55723 56389 55735 56392
rect 55677 56383 55735 56389
rect 57977 56389 57989 56392
rect 58023 56389 58035 56423
rect 57977 56383 58035 56389
rect 49513 56355 49571 56361
rect 49513 56321 49525 56355
rect 49559 56321 49571 56355
rect 55490 56352 55496 56364
rect 55451 56324 55496 56352
rect 49513 56315 49571 56321
rect 55490 56312 55496 56324
rect 55548 56312 55554 56364
rect 56870 56312 56876 56364
rect 56928 56352 56934 56364
rect 57885 56355 57943 56361
rect 57885 56352 57897 56355
rect 56928 56324 57897 56352
rect 56928 56312 56934 56324
rect 57885 56321 57897 56324
rect 57931 56321 57943 56355
rect 57885 56315 57943 56321
rect 6549 56287 6607 56293
rect 6549 56253 6561 56287
rect 6595 56284 6607 56287
rect 6914 56284 6920 56296
rect 6595 56256 6920 56284
rect 6595 56253 6607 56256
rect 6549 56247 6607 56253
rect 6914 56244 6920 56256
rect 6972 56244 6978 56296
rect 7009 56287 7067 56293
rect 7009 56253 7021 56287
rect 7055 56253 7067 56287
rect 7009 56247 7067 56253
rect 8849 56287 8907 56293
rect 8849 56253 8861 56287
rect 8895 56284 8907 56287
rect 9030 56284 9036 56296
rect 8895 56256 9036 56284
rect 8895 56253 8907 56256
rect 8849 56247 8907 56253
rect 5810 56176 5816 56228
rect 5868 56216 5874 56228
rect 7024 56216 7052 56247
rect 9030 56244 9036 56256
rect 9088 56244 9094 56296
rect 9125 56287 9183 56293
rect 9125 56253 9137 56287
rect 9171 56253 9183 56287
rect 9125 56247 9183 56253
rect 5868 56188 7052 56216
rect 5868 56176 5874 56188
rect 7098 56176 7104 56228
rect 7156 56216 7162 56228
rect 9140 56216 9168 56247
rect 13078 56244 13084 56296
rect 13136 56284 13142 56296
rect 13449 56287 13507 56293
rect 13449 56284 13461 56287
rect 13136 56256 13461 56284
rect 13136 56244 13142 56256
rect 13449 56253 13461 56256
rect 13495 56253 13507 56287
rect 13449 56247 13507 56253
rect 13538 56244 13544 56296
rect 13596 56284 13602 56296
rect 13817 56287 13875 56293
rect 13817 56284 13829 56287
rect 13596 56256 13829 56284
rect 13596 56244 13602 56256
rect 13817 56253 13829 56256
rect 13863 56253 13875 56287
rect 13817 56247 13875 56253
rect 16945 56287 17003 56293
rect 16945 56253 16957 56287
rect 16991 56284 17003 56287
rect 17126 56284 17132 56296
rect 16991 56256 17132 56284
rect 16991 56253 17003 56256
rect 16945 56247 17003 56253
rect 17126 56244 17132 56256
rect 17184 56244 17190 56296
rect 17402 56284 17408 56296
rect 17363 56256 17408 56284
rect 17402 56244 17408 56256
rect 17460 56244 17466 56296
rect 19058 56284 19064 56296
rect 19019 56256 19064 56284
rect 19058 56244 19064 56256
rect 19116 56244 19122 56296
rect 19245 56287 19303 56293
rect 19245 56253 19257 56287
rect 19291 56253 19303 56287
rect 19245 56247 19303 56253
rect 7156 56188 9168 56216
rect 7156 56176 7162 56188
rect 4706 56148 4712 56160
rect 4264 56120 4712 56148
rect 4706 56108 4712 56120
rect 4764 56148 4770 56160
rect 15102 56148 15108 56160
rect 4764 56120 15108 56148
rect 4764 56108 4770 56120
rect 15102 56108 15108 56120
rect 15160 56108 15166 56160
rect 19260 56148 19288 56247
rect 19334 56244 19340 56296
rect 19392 56284 19398 56296
rect 19521 56287 19579 56293
rect 19521 56284 19533 56287
rect 19392 56256 19533 56284
rect 19392 56244 19398 56256
rect 19521 56253 19533 56256
rect 19567 56253 19579 56287
rect 21818 56284 21824 56296
rect 21779 56256 21824 56284
rect 19521 56247 19579 56253
rect 21818 56244 21824 56256
rect 21876 56244 21882 56296
rect 23014 56284 23020 56296
rect 22975 56256 23020 56284
rect 23014 56244 23020 56256
rect 23072 56244 23078 56296
rect 26053 56287 26111 56293
rect 26053 56253 26065 56287
rect 26099 56253 26111 56287
rect 26970 56284 26976 56296
rect 26931 56256 26976 56284
rect 26053 56247 26111 56253
rect 26068 56216 26096 56247
rect 26970 56244 26976 56256
rect 27028 56244 27034 56296
rect 28350 56244 28356 56296
rect 28408 56284 28414 56296
rect 28445 56287 28503 56293
rect 28445 56284 28457 56287
rect 28408 56256 28457 56284
rect 28408 56244 28414 56256
rect 28445 56253 28457 56256
rect 28491 56253 28503 56287
rect 28445 56247 28503 56253
rect 32309 56287 32367 56293
rect 32309 56253 32321 56287
rect 32355 56284 32367 56287
rect 32398 56284 32404 56296
rect 32355 56256 32404 56284
rect 32355 56253 32367 56256
rect 32309 56247 32367 56253
rect 32398 56244 32404 56256
rect 32456 56244 32462 56296
rect 32858 56284 32864 56296
rect 32819 56256 32864 56284
rect 32858 56244 32864 56256
rect 32916 56244 32922 56296
rect 39853 56287 39911 56293
rect 39853 56253 39865 56287
rect 39899 56284 39911 56287
rect 40126 56284 40132 56296
rect 39899 56256 40132 56284
rect 39899 56253 39911 56256
rect 39853 56247 39911 56253
rect 40126 56244 40132 56256
rect 40184 56244 40190 56296
rect 40586 56284 40592 56296
rect 40547 56256 40592 56284
rect 40586 56244 40592 56256
rect 40644 56244 40650 56296
rect 42794 56284 42800 56296
rect 42755 56256 42800 56284
rect 42794 56244 42800 56256
rect 42852 56244 42858 56296
rect 49697 56287 49755 56293
rect 49697 56253 49709 56287
rect 49743 56284 49755 56287
rect 50246 56284 50252 56296
rect 49743 56256 50252 56284
rect 49743 56253 49755 56256
rect 49697 56247 49755 56253
rect 50246 56244 50252 56256
rect 50304 56244 50310 56296
rect 50341 56287 50399 56293
rect 50341 56253 50353 56287
rect 50387 56253 50399 56287
rect 56686 56284 56692 56296
rect 56647 56256 56692 56284
rect 50341 56247 50399 56253
rect 27614 56216 27620 56228
rect 26068 56188 27620 56216
rect 27614 56176 27620 56188
rect 27672 56176 27678 56228
rect 50154 56176 50160 56228
rect 50212 56216 50218 56228
rect 50356 56216 50384 56247
rect 56686 56244 56692 56256
rect 56744 56244 56750 56296
rect 50212 56188 50384 56216
rect 50212 56176 50218 56188
rect 19334 56148 19340 56160
rect 19260 56120 19340 56148
rect 19334 56108 19340 56120
rect 19392 56108 19398 56160
rect 25590 56108 25596 56160
rect 25648 56148 25654 56160
rect 26421 56151 26479 56157
rect 26421 56148 26433 56151
rect 25648 56120 26433 56148
rect 25648 56108 25654 56120
rect 26421 56117 26433 56120
rect 26467 56117 26479 56151
rect 30926 56148 30932 56160
rect 30887 56120 30932 56148
rect 26421 56111 26479 56117
rect 30926 56108 30932 56120
rect 30984 56108 30990 56160
rect 35710 56108 35716 56160
rect 35768 56148 35774 56160
rect 35989 56151 36047 56157
rect 35989 56148 36001 56151
rect 35768 56120 36001 56148
rect 35768 56108 35774 56120
rect 35989 56117 36001 56120
rect 36035 56117 36047 56151
rect 35989 56111 36047 56117
rect 46382 56108 46388 56160
rect 46440 56148 46446 56160
rect 46753 56151 46811 56157
rect 46753 56148 46765 56151
rect 46440 56120 46765 56148
rect 46440 56108 46446 56120
rect 46753 56117 46765 56120
rect 46799 56117 46811 56151
rect 46753 56111 46811 56117
rect 56226 56108 56232 56160
rect 56284 56148 56290 56160
rect 56870 56148 56876 56160
rect 56284 56120 56876 56148
rect 56284 56108 56290 56120
rect 56870 56108 56876 56120
rect 56928 56108 56934 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 6914 55904 6920 55956
rect 6972 55944 6978 55956
rect 7469 55947 7527 55953
rect 7469 55944 7481 55947
rect 6972 55916 7481 55944
rect 6972 55904 6978 55916
rect 7469 55913 7481 55916
rect 7515 55913 7527 55947
rect 9030 55944 9036 55956
rect 8991 55916 9036 55944
rect 7469 55907 7527 55913
rect 9030 55904 9036 55916
rect 9088 55904 9094 55956
rect 13078 55944 13084 55956
rect 13039 55916 13084 55944
rect 13078 55904 13084 55916
rect 13136 55904 13142 55956
rect 50246 55944 50252 55956
rect 16546 55916 50108 55944
rect 50207 55916 50252 55944
rect 9490 55836 9496 55888
rect 9548 55876 9554 55888
rect 16546 55876 16574 55916
rect 9548 55848 16574 55876
rect 9548 55836 9554 55848
rect 19058 55836 19064 55888
rect 19116 55876 19122 55888
rect 19429 55879 19487 55885
rect 19429 55876 19441 55879
rect 19116 55848 19441 55876
rect 19116 55836 19122 55848
rect 19429 55845 19441 55848
rect 19475 55845 19487 55879
rect 20438 55876 20444 55888
rect 20399 55848 20444 55876
rect 19429 55839 19487 55845
rect 20438 55836 20444 55848
rect 20496 55836 20502 55888
rect 28166 55836 28172 55888
rect 28224 55876 28230 55888
rect 32398 55876 32404 55888
rect 28224 55848 30604 55876
rect 32359 55848 32404 55876
rect 28224 55836 28230 55848
rect 9508 55808 9536 55836
rect 2608 55780 6914 55808
rect 1486 55740 1492 55752
rect 1447 55712 1492 55740
rect 1486 55700 1492 55712
rect 1544 55700 1550 55752
rect 2608 55749 2636 55780
rect 2593 55743 2651 55749
rect 2593 55709 2605 55743
rect 2639 55709 2651 55743
rect 2593 55703 2651 55709
rect 3694 55700 3700 55752
rect 3752 55740 3758 55752
rect 3789 55743 3847 55749
rect 3789 55740 3801 55743
rect 3752 55712 3801 55740
rect 3752 55700 3758 55712
rect 3789 55709 3801 55712
rect 3835 55709 3847 55743
rect 3789 55703 3847 55709
rect 2038 55672 2044 55684
rect 1999 55644 2044 55672
rect 2038 55632 2044 55644
rect 2096 55632 2102 55684
rect 2685 55675 2743 55681
rect 2685 55641 2697 55675
rect 2731 55672 2743 55675
rect 3973 55675 4031 55681
rect 3973 55672 3985 55675
rect 2731 55644 3985 55672
rect 2731 55641 2743 55644
rect 2685 55635 2743 55641
rect 3973 55641 3985 55644
rect 4019 55641 4031 55675
rect 5629 55675 5687 55681
rect 5629 55672 5641 55675
rect 3973 55635 4031 55641
rect 5460 55644 5641 55672
rect 2590 55564 2596 55616
rect 2648 55604 2654 55616
rect 5460 55604 5488 55644
rect 5629 55641 5641 55644
rect 5675 55641 5687 55675
rect 5629 55635 5687 55641
rect 2648 55576 5488 55604
rect 6886 55604 6914 55780
rect 7392 55780 9536 55808
rect 15749 55811 15807 55817
rect 7392 55749 7420 55780
rect 15749 55777 15761 55811
rect 15795 55808 15807 55811
rect 16022 55808 16028 55820
rect 15795 55780 16028 55808
rect 15795 55777 15807 55780
rect 15749 55771 15807 55777
rect 16022 55768 16028 55780
rect 16080 55768 16086 55820
rect 16114 55768 16120 55820
rect 16172 55808 16178 55820
rect 16209 55811 16267 55817
rect 16209 55808 16221 55811
rect 16172 55780 16221 55808
rect 16172 55768 16178 55780
rect 16209 55777 16221 55780
rect 16255 55777 16267 55811
rect 20456 55808 20484 55836
rect 20456 55780 21036 55808
rect 16209 55771 16267 55777
rect 7377 55743 7435 55749
rect 7377 55709 7389 55743
rect 7423 55709 7435 55743
rect 8938 55740 8944 55752
rect 8899 55712 8944 55740
rect 7377 55703 7435 55709
rect 8938 55700 8944 55712
rect 8996 55700 9002 55752
rect 12986 55740 12992 55752
rect 12947 55712 12992 55740
rect 12986 55700 12992 55712
rect 13044 55700 13050 55752
rect 15102 55740 15108 55752
rect 15063 55712 15108 55740
rect 15102 55700 15108 55712
rect 15160 55700 15166 55752
rect 21008 55749 21036 55780
rect 21928 55780 22968 55808
rect 20901 55743 20959 55749
rect 20901 55709 20913 55743
rect 20947 55709 20959 55743
rect 20901 55703 20959 55709
rect 20993 55743 21051 55749
rect 20993 55709 21005 55743
rect 21039 55709 21051 55743
rect 21818 55740 21824 55752
rect 20993 55703 21051 55709
rect 21100 55712 21824 55740
rect 15197 55675 15255 55681
rect 15197 55641 15209 55675
rect 15243 55672 15255 55675
rect 15933 55675 15991 55681
rect 15933 55672 15945 55675
rect 15243 55644 15945 55672
rect 15243 55641 15255 55644
rect 15197 55635 15255 55641
rect 15933 55641 15945 55644
rect 15979 55641 15991 55675
rect 20916 55672 20944 55703
rect 21100 55672 21128 55712
rect 21818 55700 21824 55712
rect 21876 55700 21882 55752
rect 21928 55749 21956 55780
rect 21913 55743 21971 55749
rect 21913 55709 21925 55743
rect 21959 55709 21971 55743
rect 21913 55703 21971 55709
rect 22741 55743 22799 55749
rect 22741 55709 22753 55743
rect 22787 55709 22799 55743
rect 22741 55703 22799 55709
rect 20916 55644 21128 55672
rect 21177 55675 21235 55681
rect 15933 55635 15991 55641
rect 21177 55641 21189 55675
rect 21223 55672 21235 55675
rect 22756 55672 22784 55703
rect 21223 55644 22784 55672
rect 21223 55641 21235 55644
rect 21177 55635 21235 55641
rect 16574 55604 16580 55616
rect 6886 55576 16580 55604
rect 2648 55564 2654 55576
rect 16574 55564 16580 55576
rect 16632 55604 16638 55616
rect 17310 55604 17316 55616
rect 16632 55576 17316 55604
rect 16632 55564 16638 55576
rect 17310 55564 17316 55576
rect 17368 55564 17374 55616
rect 21266 55564 21272 55616
rect 21324 55604 21330 55616
rect 22097 55607 22155 55613
rect 22097 55604 22109 55607
rect 21324 55576 22109 55604
rect 21324 55564 21330 55576
rect 22097 55573 22109 55576
rect 22143 55573 22155 55607
rect 22554 55604 22560 55616
rect 22515 55576 22560 55604
rect 22097 55567 22155 55573
rect 22554 55564 22560 55576
rect 22612 55564 22618 55616
rect 22940 55604 22968 55780
rect 23014 55768 23020 55820
rect 23072 55808 23078 55820
rect 24949 55811 25007 55817
rect 24949 55808 24961 55811
rect 23072 55780 24961 55808
rect 23072 55768 23078 55780
rect 24949 55777 24961 55780
rect 24995 55808 25007 55811
rect 30009 55811 30067 55817
rect 24995 55780 25084 55808
rect 24995 55777 25007 55780
rect 24949 55771 25007 55777
rect 25056 55752 25084 55780
rect 30009 55777 30021 55811
rect 30055 55808 30067 55811
rect 30190 55808 30196 55820
rect 30055 55780 30196 55808
rect 30055 55777 30067 55780
rect 30009 55771 30067 55777
rect 30190 55768 30196 55780
rect 30248 55768 30254 55820
rect 30282 55768 30288 55820
rect 30340 55808 30346 55820
rect 30469 55811 30527 55817
rect 30469 55808 30481 55811
rect 30340 55780 30481 55808
rect 30340 55768 30346 55780
rect 30469 55777 30481 55780
rect 30515 55777 30527 55811
rect 30576 55808 30604 55848
rect 32398 55836 32404 55848
rect 32456 55836 32462 55888
rect 35161 55879 35219 55885
rect 35161 55845 35173 55879
rect 35207 55876 35219 55879
rect 35802 55876 35808 55888
rect 35207 55848 35808 55876
rect 35207 55845 35219 55848
rect 35161 55839 35219 55845
rect 35802 55836 35808 55848
rect 35860 55836 35866 55888
rect 40126 55876 40132 55888
rect 40087 55848 40132 55876
rect 40126 55836 40132 55848
rect 40184 55836 40190 55888
rect 50080 55876 50108 55916
rect 50246 55904 50252 55916
rect 50304 55904 50310 55956
rect 55398 55904 55404 55956
rect 55456 55944 55462 55956
rect 57238 55944 57244 55956
rect 55456 55916 57244 55944
rect 55456 55904 55462 55916
rect 57238 55904 57244 55916
rect 57296 55904 57302 55956
rect 56226 55876 56232 55888
rect 40512 55848 45554 55876
rect 50080 55848 56232 55876
rect 40512 55808 40540 55848
rect 30576 55780 40540 55808
rect 30469 55771 30527 55777
rect 42242 55768 42248 55820
rect 42300 55808 42306 55820
rect 42429 55811 42487 55817
rect 42429 55808 42441 55811
rect 42300 55780 42441 55808
rect 42300 55768 42306 55780
rect 42429 55777 42441 55780
rect 42475 55777 42487 55811
rect 43806 55808 43812 55820
rect 43767 55780 43812 55808
rect 42429 55771 42487 55777
rect 43806 55768 43812 55780
rect 43864 55768 43870 55820
rect 25038 55700 25044 55752
rect 25096 55740 25102 55752
rect 27065 55743 27123 55749
rect 27065 55740 27077 55743
rect 25096 55712 27077 55740
rect 25096 55700 25102 55712
rect 27065 55709 27077 55712
rect 27111 55709 27123 55743
rect 27065 55703 27123 55709
rect 27154 55700 27160 55752
rect 27212 55740 27218 55752
rect 27321 55743 27379 55749
rect 27321 55740 27333 55743
rect 27212 55712 27333 55740
rect 27212 55700 27218 55712
rect 27321 55709 27333 55712
rect 27367 55709 27379 55743
rect 27321 55703 27379 55709
rect 32214 55700 32220 55752
rect 32272 55740 32278 55752
rect 32309 55743 32367 55749
rect 32309 55740 32321 55743
rect 32272 55712 32321 55740
rect 32272 55700 32278 55712
rect 32309 55709 32321 55712
rect 32355 55740 32367 55743
rect 33137 55743 33195 55749
rect 33137 55740 33149 55743
rect 32355 55712 33149 55740
rect 32355 55709 32367 55712
rect 32309 55703 32367 55709
rect 33137 55709 33149 55712
rect 33183 55709 33195 55743
rect 33137 55703 33195 55709
rect 35069 55743 35127 55749
rect 35069 55709 35081 55743
rect 35115 55740 35127 55743
rect 35342 55740 35348 55752
rect 35115 55712 35348 55740
rect 35115 55709 35127 55712
rect 35069 55703 35127 55709
rect 35342 55700 35348 55712
rect 35400 55700 35406 55752
rect 35710 55740 35716 55752
rect 35671 55712 35716 55740
rect 35710 55700 35716 55712
rect 35768 55700 35774 55752
rect 40034 55740 40040 55752
rect 39995 55712 40040 55740
rect 40034 55700 40040 55712
rect 40092 55700 40098 55752
rect 25216 55675 25274 55681
rect 25216 55641 25228 55675
rect 25262 55672 25274 55675
rect 25406 55672 25412 55684
rect 25262 55644 25412 55672
rect 25262 55641 25274 55644
rect 25216 55635 25274 55641
rect 25406 55632 25412 55644
rect 25464 55632 25470 55684
rect 30193 55675 30251 55681
rect 26206 55644 28580 55672
rect 26206 55604 26234 55644
rect 26326 55604 26332 55616
rect 22940 55576 26234 55604
rect 26287 55576 26332 55604
rect 26326 55564 26332 55576
rect 26384 55564 26390 55616
rect 28442 55604 28448 55616
rect 28403 55576 28448 55604
rect 28442 55564 28448 55576
rect 28500 55564 28506 55616
rect 28552 55604 28580 55644
rect 30193 55641 30205 55675
rect 30239 55672 30251 55675
rect 30926 55672 30932 55684
rect 30239 55644 30932 55672
rect 30239 55641 30251 55644
rect 30193 55635 30251 55641
rect 30926 55632 30932 55644
rect 30984 55632 30990 55684
rect 33229 55675 33287 55681
rect 33229 55641 33241 55675
rect 33275 55672 33287 55675
rect 35897 55675 35955 55681
rect 33275 55644 35296 55672
rect 33275 55641 33287 55644
rect 33229 55635 33287 55641
rect 33594 55604 33600 55616
rect 28552 55576 33600 55604
rect 33594 55564 33600 55576
rect 33652 55564 33658 55616
rect 35268 55604 35296 55644
rect 35897 55641 35909 55675
rect 35943 55672 35955 55675
rect 36262 55672 36268 55684
rect 35943 55644 36268 55672
rect 35943 55641 35955 55644
rect 35897 55635 35955 55641
rect 36262 55632 36268 55644
rect 36320 55632 36326 55684
rect 36722 55632 36728 55684
rect 36780 55672 36786 55684
rect 37553 55675 37611 55681
rect 37553 55672 37565 55675
rect 36780 55644 37565 55672
rect 36780 55632 36786 55644
rect 37553 55641 37565 55644
rect 37599 55641 37611 55675
rect 42610 55672 42616 55684
rect 42571 55644 42616 55672
rect 37553 55635 37611 55641
rect 42610 55632 42616 55644
rect 42668 55632 42674 55684
rect 42794 55604 42800 55616
rect 35268 55576 42800 55604
rect 42794 55564 42800 55576
rect 42852 55564 42858 55616
rect 45526 55604 45554 55848
rect 56226 55836 56232 55848
rect 56284 55836 56290 55888
rect 57422 55876 57428 55888
rect 56336 55848 57428 55876
rect 46198 55808 46204 55820
rect 46159 55780 46204 55808
rect 46198 55768 46204 55780
rect 46256 55768 46262 55820
rect 46382 55808 46388 55820
rect 46343 55780 46388 55808
rect 46382 55768 46388 55780
rect 46440 55768 46446 55820
rect 47026 55808 47032 55820
rect 46987 55780 47032 55808
rect 47026 55768 47032 55780
rect 47084 55768 47090 55820
rect 54757 55811 54815 55817
rect 54757 55777 54769 55811
rect 54803 55808 54815 55811
rect 56042 55808 56048 55820
rect 54803 55780 56048 55808
rect 54803 55777 54815 55780
rect 54757 55771 54815 55777
rect 56042 55768 56048 55780
rect 56100 55768 56106 55820
rect 56336 55817 56364 55848
rect 57422 55836 57428 55848
rect 57480 55836 57486 55888
rect 56321 55811 56379 55817
rect 56321 55777 56333 55811
rect 56367 55777 56379 55811
rect 56321 55771 56379 55777
rect 56502 55768 56508 55820
rect 56560 55808 56566 55820
rect 56781 55811 56839 55817
rect 56781 55808 56793 55811
rect 56560 55780 56793 55808
rect 56560 55768 56566 55780
rect 56781 55777 56793 55780
rect 56827 55777 56839 55811
rect 56781 55771 56839 55777
rect 47854 55700 47860 55752
rect 47912 55740 47918 55752
rect 50157 55743 50215 55749
rect 50157 55740 50169 55743
rect 47912 55712 50169 55740
rect 47912 55700 47918 55712
rect 50157 55709 50169 55712
rect 50203 55709 50215 55743
rect 52914 55740 52920 55752
rect 52875 55712 52920 55740
rect 50157 55703 50215 55709
rect 52914 55700 52920 55712
rect 52972 55700 52978 55752
rect 55306 55700 55312 55752
rect 55364 55740 55370 55752
rect 55674 55740 55680 55752
rect 55364 55712 55680 55740
rect 55364 55700 55370 55712
rect 55674 55700 55680 55712
rect 55732 55700 55738 55752
rect 53101 55675 53159 55681
rect 53101 55641 53113 55675
rect 53147 55672 53159 55675
rect 54662 55672 54668 55684
rect 53147 55644 54668 55672
rect 53147 55641 53159 55644
rect 53101 55635 53159 55641
rect 54662 55632 54668 55644
rect 54720 55632 54726 55684
rect 55769 55675 55827 55681
rect 55769 55641 55781 55675
rect 55815 55672 55827 55675
rect 56505 55675 56563 55681
rect 56505 55672 56517 55675
rect 55815 55644 56517 55672
rect 55815 55641 55827 55644
rect 55769 55635 55827 55641
rect 56505 55641 56517 55644
rect 56551 55641 56563 55675
rect 56505 55635 56563 55641
rect 56778 55604 56784 55616
rect 45526 55576 56784 55604
rect 56778 55564 56784 55576
rect 56836 55564 56842 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 21818 55360 21824 55412
rect 21876 55400 21882 55412
rect 23201 55403 23259 55409
rect 21876 55372 22692 55400
rect 21876 55360 21882 55372
rect 2866 55332 2872 55344
rect 2332 55304 2872 55332
rect 2332 55273 2360 55304
rect 2866 55292 2872 55304
rect 2924 55292 2930 55344
rect 17954 55332 17960 55344
rect 17696 55304 17960 55332
rect 17696 55273 17724 55304
rect 17954 55292 17960 55304
rect 18012 55292 18018 55344
rect 22088 55335 22146 55341
rect 22088 55301 22100 55335
rect 22134 55332 22146 55335
rect 22554 55332 22560 55344
rect 22134 55304 22560 55332
rect 22134 55301 22146 55304
rect 22088 55295 22146 55301
rect 22554 55292 22560 55304
rect 22612 55292 22618 55344
rect 22664 55332 22692 55372
rect 23201 55369 23213 55403
rect 23247 55400 23259 55403
rect 23658 55400 23664 55412
rect 23247 55372 23664 55400
rect 23247 55369 23259 55372
rect 23201 55363 23259 55369
rect 23658 55360 23664 55372
rect 23716 55360 23722 55412
rect 25406 55400 25412 55412
rect 25367 55372 25412 55400
rect 25406 55360 25412 55372
rect 25464 55360 25470 55412
rect 26421 55403 26479 55409
rect 26421 55369 26433 55403
rect 26467 55400 26479 55403
rect 36262 55400 36268 55412
rect 26467 55372 29500 55400
rect 36223 55372 36268 55400
rect 26467 55369 26479 55372
rect 26421 55363 26479 55369
rect 27338 55332 27344 55344
rect 22664 55304 27344 55332
rect 27338 55292 27344 55304
rect 27396 55292 27402 55344
rect 28534 55332 28540 55344
rect 27448 55304 28540 55332
rect 2317 55267 2375 55273
rect 2317 55233 2329 55267
rect 2363 55233 2375 55267
rect 2317 55227 2375 55233
rect 17681 55267 17739 55273
rect 17681 55233 17693 55267
rect 17727 55233 17739 55267
rect 21266 55264 21272 55276
rect 21227 55236 21272 55264
rect 17681 55227 17739 55233
rect 21266 55224 21272 55236
rect 21324 55224 21330 55276
rect 21821 55267 21879 55273
rect 21821 55233 21833 55267
rect 21867 55264 21879 55267
rect 21910 55264 21916 55276
rect 21867 55236 21916 55264
rect 21867 55233 21879 55236
rect 21821 55227 21879 55233
rect 21910 55224 21916 55236
rect 21968 55224 21974 55276
rect 25590 55264 25596 55276
rect 25551 55236 25596 55264
rect 25590 55224 25596 55236
rect 25648 55224 25654 55276
rect 26142 55224 26148 55276
rect 26200 55264 26206 55276
rect 27448 55273 27476 55304
rect 28534 55292 28540 55304
rect 28592 55292 28598 55344
rect 26237 55267 26295 55273
rect 26237 55264 26249 55267
rect 26200 55236 26249 55264
rect 26200 55224 26206 55236
rect 26237 55233 26249 55236
rect 26283 55233 26295 55267
rect 26237 55227 26295 55233
rect 27433 55267 27491 55273
rect 27433 55233 27445 55267
rect 27479 55233 27491 55267
rect 27433 55227 27491 55233
rect 27700 55267 27758 55273
rect 27700 55233 27712 55267
rect 27746 55264 27758 55267
rect 29270 55264 29276 55276
rect 27746 55236 29276 55264
rect 27746 55233 27758 55236
rect 27700 55227 27758 55233
rect 29270 55224 29276 55236
rect 29328 55224 29334 55276
rect 29472 55273 29500 55372
rect 36262 55360 36268 55372
rect 36320 55360 36326 55412
rect 40034 55360 40040 55412
rect 40092 55400 40098 55412
rect 54662 55400 54668 55412
rect 40092 55372 45554 55400
rect 54623 55372 54668 55400
rect 40092 55360 40098 55372
rect 45526 55332 45554 55372
rect 54662 55360 54668 55372
rect 54720 55360 54726 55412
rect 56594 55400 56600 55412
rect 55508 55372 56600 55400
rect 55306 55332 55312 55344
rect 45526 55304 55312 55332
rect 55306 55292 55312 55304
rect 55364 55292 55370 55344
rect 29457 55267 29515 55273
rect 29457 55233 29469 55267
rect 29503 55233 29515 55267
rect 36170 55264 36176 55276
rect 36131 55236 36176 55264
rect 29457 55227 29515 55233
rect 36170 55224 36176 55236
rect 36228 55224 36234 55276
rect 54573 55267 54631 55273
rect 54573 55233 54585 55267
rect 54619 55264 54631 55267
rect 54619 55236 55352 55264
rect 54619 55233 54631 55236
rect 54573 55227 54631 55233
rect 2501 55199 2559 55205
rect 2501 55165 2513 55199
rect 2547 55196 2559 55199
rect 3786 55196 3792 55208
rect 2547 55168 3792 55196
rect 2547 55165 2559 55168
rect 2501 55159 2559 55165
rect 3786 55156 3792 55168
rect 3844 55156 3850 55208
rect 3970 55196 3976 55208
rect 3931 55168 3976 55196
rect 3970 55156 3976 55168
rect 4028 55156 4034 55208
rect 17862 55196 17868 55208
rect 17823 55168 17868 55196
rect 17862 55156 17868 55168
rect 17920 55156 17926 55208
rect 19242 55196 19248 55208
rect 19203 55168 19248 55196
rect 19242 55156 19248 55168
rect 19300 55156 19306 55208
rect 26050 55196 26056 55208
rect 26011 55168 26056 55196
rect 26050 55156 26056 55168
rect 26108 55156 26114 55208
rect 28534 55156 28540 55208
rect 28592 55196 28598 55208
rect 29546 55196 29552 55208
rect 28592 55168 29552 55196
rect 28592 55156 28598 55168
rect 29546 55156 29552 55168
rect 29604 55156 29610 55208
rect 29270 55128 29276 55140
rect 29231 55100 29276 55128
rect 29270 55088 29276 55100
rect 29328 55088 29334 55140
rect 55324 55128 55352 55236
rect 55398 55224 55404 55276
rect 55456 55224 55462 55276
rect 55508 55273 55536 55372
rect 56594 55360 56600 55372
rect 56652 55360 56658 55412
rect 56778 55360 56784 55412
rect 56836 55400 56842 55412
rect 57974 55400 57980 55412
rect 56836 55372 57468 55400
rect 57935 55372 57980 55400
rect 56836 55360 56842 55372
rect 57330 55332 57336 55344
rect 57291 55304 57336 55332
rect 57330 55292 57336 55304
rect 57388 55292 57394 55344
rect 55493 55267 55551 55273
rect 55493 55233 55505 55267
rect 55539 55233 55551 55267
rect 57440 55264 57468 55372
rect 57974 55360 57980 55372
rect 58032 55360 58038 55412
rect 57885 55267 57943 55273
rect 57885 55264 57897 55267
rect 57440 55236 57897 55264
rect 55493 55227 55551 55233
rect 57885 55233 57897 55236
rect 57931 55233 57943 55267
rect 57885 55227 57943 55233
rect 55416 55196 55444 55224
rect 55677 55199 55735 55205
rect 55677 55196 55689 55199
rect 55416 55168 55689 55196
rect 55677 55165 55689 55168
rect 55723 55165 55735 55199
rect 55677 55159 55735 55165
rect 56594 55128 56600 55140
rect 55324 55100 56600 55128
rect 56594 55088 56600 55100
rect 56652 55088 56658 55140
rect 21082 55060 21088 55072
rect 21043 55032 21088 55060
rect 21082 55020 21088 55032
rect 21140 55020 21146 55072
rect 27614 55020 27620 55072
rect 27672 55060 27678 55072
rect 28074 55060 28080 55072
rect 27672 55032 28080 55060
rect 27672 55020 27678 55032
rect 28074 55020 28080 55032
rect 28132 55060 28138 55072
rect 28813 55063 28871 55069
rect 28813 55060 28825 55063
rect 28132 55032 28825 55060
rect 28132 55020 28138 55032
rect 28813 55029 28825 55032
rect 28859 55029 28871 55063
rect 28813 55023 28871 55029
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 2130 54816 2136 54868
rect 2188 54856 2194 54868
rect 2593 54859 2651 54865
rect 2593 54856 2605 54859
rect 2188 54828 2605 54856
rect 2188 54816 2194 54828
rect 2593 54825 2605 54828
rect 2639 54825 2651 54859
rect 2593 54819 2651 54825
rect 3786 54816 3792 54868
rect 3844 54856 3850 54868
rect 3881 54859 3939 54865
rect 3881 54856 3893 54859
rect 3844 54828 3893 54856
rect 3844 54816 3850 54828
rect 3881 54825 3893 54828
rect 3927 54825 3939 54859
rect 19334 54856 19340 54868
rect 19295 54828 19340 54856
rect 3881 54819 3939 54825
rect 19334 54816 19340 54828
rect 19392 54816 19398 54868
rect 27433 54859 27491 54865
rect 27433 54825 27445 54859
rect 27479 54856 27491 54859
rect 27614 54856 27620 54868
rect 27479 54828 27620 54856
rect 27479 54825 27491 54828
rect 27433 54819 27491 54825
rect 27614 54816 27620 54828
rect 27672 54816 27678 54868
rect 27890 54816 27896 54868
rect 27948 54856 27954 54868
rect 28353 54859 28411 54865
rect 28353 54856 28365 54859
rect 27948 54828 28365 54856
rect 27948 54816 27954 54828
rect 28353 54825 28365 54828
rect 28399 54856 28411 54859
rect 28442 54856 28448 54868
rect 28399 54828 28448 54856
rect 28399 54825 28411 54828
rect 28353 54819 28411 54825
rect 28442 54816 28448 54828
rect 28500 54816 28506 54868
rect 26050 54680 26056 54732
rect 26108 54720 26114 54732
rect 28169 54723 28227 54729
rect 28169 54720 28181 54723
rect 26108 54692 28181 54720
rect 26108 54680 26114 54692
rect 28169 54689 28181 54692
rect 28215 54720 28227 54723
rect 28994 54720 29000 54732
rect 28215 54692 29000 54720
rect 28215 54689 28227 54692
rect 28169 54683 28227 54689
rect 28994 54680 29000 54692
rect 29052 54680 29058 54732
rect 58158 54720 58164 54732
rect 58119 54692 58164 54720
rect 58158 54680 58164 54692
rect 58216 54680 58222 54732
rect 2501 54655 2559 54661
rect 2501 54621 2513 54655
rect 2547 54652 2559 54655
rect 3326 54652 3332 54664
rect 2547 54624 3332 54652
rect 2547 54621 2559 54624
rect 2501 54615 2559 54621
rect 3326 54612 3332 54624
rect 3384 54612 3390 54664
rect 3789 54655 3847 54661
rect 3789 54621 3801 54655
rect 3835 54652 3847 54655
rect 3970 54652 3976 54664
rect 3835 54624 3976 54652
rect 3835 54621 3847 54624
rect 3789 54615 3847 54621
rect 3970 54612 3976 54624
rect 4028 54612 4034 54664
rect 19150 54612 19156 54664
rect 19208 54652 19214 54664
rect 19245 54655 19303 54661
rect 19245 54652 19257 54655
rect 19208 54624 19257 54652
rect 19208 54612 19214 54624
rect 19245 54621 19257 54624
rect 19291 54621 19303 54655
rect 19245 54615 19303 54621
rect 20073 54655 20131 54661
rect 20073 54621 20085 54655
rect 20119 54652 20131 54655
rect 21910 54652 21916 54664
rect 20119 54624 21916 54652
rect 20119 54621 20131 54624
rect 20073 54615 20131 54621
rect 21910 54612 21916 54624
rect 21968 54612 21974 54664
rect 28353 54655 28411 54661
rect 28353 54652 28365 54655
rect 27264 54624 28365 54652
rect 20340 54587 20398 54593
rect 20340 54553 20352 54587
rect 20386 54584 20398 54587
rect 21082 54584 21088 54596
rect 20386 54556 21088 54584
rect 20386 54553 20398 54556
rect 20340 54547 20398 54553
rect 21082 54544 21088 54556
rect 21140 54544 21146 54596
rect 26970 54544 26976 54596
rect 27028 54584 27034 54596
rect 27264 54593 27292 54624
rect 28353 54621 28365 54624
rect 28399 54621 28411 54655
rect 29546 54652 29552 54664
rect 29507 54624 29552 54652
rect 28353 54615 28411 54621
rect 29546 54612 29552 54624
rect 29604 54612 29610 54664
rect 56318 54652 56324 54664
rect 56279 54624 56324 54652
rect 56318 54612 56324 54624
rect 56376 54612 56382 54664
rect 27249 54587 27307 54593
rect 27249 54584 27261 54587
rect 27028 54556 27261 54584
rect 27028 54544 27034 54556
rect 27249 54553 27261 54556
rect 27295 54553 27307 54587
rect 28074 54584 28080 54596
rect 28035 54556 28080 54584
rect 27249 54547 27307 54553
rect 28074 54544 28080 54556
rect 28132 54544 28138 54596
rect 29638 54544 29644 54596
rect 29696 54584 29702 54596
rect 29794 54587 29852 54593
rect 29794 54584 29806 54587
rect 29696 54556 29806 54584
rect 29696 54544 29702 54556
rect 29794 54553 29806 54556
rect 29840 54553 29852 54587
rect 29794 54547 29852 54553
rect 33229 54587 33287 54593
rect 33229 54553 33241 54587
rect 33275 54584 33287 54587
rect 34422 54584 34428 54596
rect 33275 54556 34428 54584
rect 33275 54553 33287 54556
rect 33229 54547 33287 54553
rect 34422 54544 34428 54556
rect 34480 54544 34486 54596
rect 56505 54587 56563 54593
rect 56505 54553 56517 54587
rect 56551 54584 56563 54587
rect 56962 54584 56968 54596
rect 56551 54556 56968 54584
rect 56551 54553 56563 54556
rect 56505 54547 56563 54553
rect 56962 54544 56968 54556
rect 57020 54544 57026 54596
rect 19978 54476 19984 54528
rect 20036 54516 20042 54528
rect 21453 54519 21511 54525
rect 21453 54516 21465 54519
rect 20036 54488 21465 54516
rect 20036 54476 20042 54488
rect 21453 54485 21465 54488
rect 21499 54485 21511 54519
rect 21453 54479 21511 54485
rect 27430 54476 27436 54528
rect 27488 54525 27494 54528
rect 27488 54519 27507 54525
rect 27495 54485 27507 54519
rect 27488 54479 27507 54485
rect 27617 54519 27675 54525
rect 27617 54485 27629 54519
rect 27663 54516 27675 54519
rect 28442 54516 28448 54528
rect 27663 54488 28448 54516
rect 27663 54485 27675 54488
rect 27617 54479 27675 54485
rect 27488 54476 27494 54479
rect 28442 54476 28448 54488
rect 28500 54476 28506 54528
rect 28537 54519 28595 54525
rect 28537 54485 28549 54519
rect 28583 54516 28595 54519
rect 28718 54516 28724 54528
rect 28583 54488 28724 54516
rect 28583 54485 28595 54488
rect 28537 54479 28595 54485
rect 28718 54476 28724 54488
rect 28776 54476 28782 54528
rect 28994 54476 29000 54528
rect 29052 54516 29058 54528
rect 30929 54519 30987 54525
rect 30929 54516 30941 54519
rect 29052 54488 30941 54516
rect 29052 54476 29058 54488
rect 30929 54485 30941 54488
rect 30975 54485 30987 54519
rect 30929 54479 30987 54485
rect 33321 54519 33379 54525
rect 33321 54485 33333 54519
rect 33367 54516 33379 54519
rect 52914 54516 52920 54528
rect 33367 54488 52920 54516
rect 33367 54485 33379 54488
rect 33321 54479 33379 54485
rect 52914 54476 52920 54488
rect 52972 54476 52978 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 29638 54312 29644 54324
rect 29599 54284 29644 54312
rect 29638 54272 29644 54284
rect 29696 54272 29702 54324
rect 56962 54312 56968 54324
rect 56923 54284 56968 54312
rect 56962 54272 56968 54284
rect 57020 54272 57026 54324
rect 26326 54244 26332 54256
rect 25976 54216 26332 54244
rect 25976 54185 26004 54216
rect 26326 54204 26332 54216
rect 26384 54204 26390 54256
rect 29178 54244 29184 54256
rect 28000 54216 29184 54244
rect 25961 54179 26019 54185
rect 25961 54145 25973 54179
rect 26007 54145 26019 54179
rect 25961 54139 26019 54145
rect 26053 54179 26111 54185
rect 26053 54145 26065 54179
rect 26099 54176 26111 54179
rect 26142 54176 26148 54188
rect 26099 54148 26148 54176
rect 26099 54145 26111 54148
rect 26053 54139 26111 54145
rect 26142 54136 26148 54148
rect 26200 54136 26206 54188
rect 27890 54176 27896 54188
rect 27851 54148 27896 54176
rect 27890 54136 27896 54148
rect 27948 54136 27954 54188
rect 28000 54185 28028 54216
rect 29178 54204 29184 54216
rect 29236 54204 29242 54256
rect 27985 54179 28043 54185
rect 27985 54145 27997 54179
rect 28031 54145 28043 54179
rect 27985 54139 28043 54145
rect 28442 54136 28448 54188
rect 28500 54176 28506 54188
rect 28813 54179 28871 54185
rect 28813 54176 28825 54179
rect 28500 54148 28825 54176
rect 28500 54136 28506 54148
rect 28813 54145 28825 54148
rect 28859 54145 28871 54179
rect 28813 54139 28871 54145
rect 28905 54179 28963 54185
rect 28905 54145 28917 54179
rect 28951 54176 28963 54179
rect 29656 54176 29684 54272
rect 56318 54204 56324 54256
rect 56376 54244 56382 54256
rect 56376 54216 58112 54244
rect 56376 54204 56382 54216
rect 28951 54148 29684 54176
rect 29825 54179 29883 54185
rect 28951 54145 28963 54148
rect 28905 54139 28963 54145
rect 29825 54145 29837 54179
rect 29871 54145 29883 54179
rect 56226 54176 56232 54188
rect 56187 54148 56232 54176
rect 29825 54139 29883 54145
rect 28994 54108 29000 54120
rect 28955 54080 29000 54108
rect 28994 54068 29000 54080
rect 29052 54068 29058 54120
rect 29086 54068 29092 54120
rect 29144 54108 29150 54120
rect 29144 54080 29189 54108
rect 29144 54068 29150 54080
rect 28169 54043 28227 54049
rect 28169 54009 28181 54043
rect 28215 54040 28227 54043
rect 29840 54040 29868 54139
rect 56226 54136 56232 54148
rect 56284 54136 56290 54188
rect 56870 54176 56876 54188
rect 56831 54148 56876 54176
rect 56870 54136 56876 54148
rect 56928 54136 56934 54188
rect 58084 54185 58112 54216
rect 58069 54179 58127 54185
rect 58069 54145 58081 54179
rect 58115 54145 58127 54179
rect 58069 54139 58127 54145
rect 28215 54012 29868 54040
rect 28215 54009 28227 54012
rect 28169 54003 28227 54009
rect 26234 53932 26240 53984
rect 26292 53972 26298 53984
rect 28629 53975 28687 53981
rect 26292 53944 26337 53972
rect 26292 53932 26298 53944
rect 28629 53941 28641 53975
rect 28675 53972 28687 53975
rect 29638 53972 29644 53984
rect 28675 53944 29644 53972
rect 28675 53941 28687 53944
rect 28629 53935 28687 53941
rect 29638 53932 29644 53944
rect 29696 53932 29702 53984
rect 56321 53975 56379 53981
rect 56321 53941 56333 53975
rect 56367 53972 56379 53975
rect 56502 53972 56508 53984
rect 56367 53944 56508 53972
rect 56367 53941 56379 53944
rect 56321 53935 56379 53941
rect 56502 53932 56508 53944
rect 56560 53932 56566 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 27430 53728 27436 53780
rect 27488 53768 27494 53780
rect 27525 53771 27583 53777
rect 27525 53768 27537 53771
rect 27488 53740 27537 53768
rect 27488 53728 27494 53740
rect 27525 53737 27537 53740
rect 27571 53737 27583 53771
rect 27525 53731 27583 53737
rect 28353 53771 28411 53777
rect 28353 53737 28365 53771
rect 28399 53768 28411 53771
rect 29086 53768 29092 53780
rect 28399 53740 29092 53768
rect 28399 53737 28411 53740
rect 28353 53731 28411 53737
rect 29086 53728 29092 53740
rect 29144 53728 29150 53780
rect 26326 53660 26332 53712
rect 26384 53700 26390 53712
rect 26973 53703 27031 53709
rect 26973 53700 26985 53703
rect 26384 53672 26985 53700
rect 26384 53660 26390 53672
rect 26973 53669 26985 53672
rect 27019 53700 27031 53703
rect 27246 53700 27252 53712
rect 27019 53672 27252 53700
rect 27019 53669 27031 53672
rect 26973 53663 27031 53669
rect 27246 53660 27252 53672
rect 27304 53660 27310 53712
rect 25038 53592 25044 53644
rect 25096 53632 25102 53644
rect 25133 53635 25191 53641
rect 25133 53632 25145 53635
rect 25096 53604 25145 53632
rect 25096 53592 25102 53604
rect 25133 53601 25145 53604
rect 25179 53601 25191 53635
rect 56502 53632 56508 53644
rect 56463 53604 56508 53632
rect 25133 53595 25191 53601
rect 56502 53592 56508 53604
rect 56560 53592 56566 53644
rect 58158 53632 58164 53644
rect 58119 53604 58164 53632
rect 58158 53592 58164 53604
rect 58216 53592 58222 53644
rect 1946 53524 1952 53576
rect 2004 53564 2010 53576
rect 2225 53567 2283 53573
rect 2225 53564 2237 53567
rect 2004 53536 2237 53564
rect 2004 53524 2010 53536
rect 2225 53533 2237 53536
rect 2271 53533 2283 53567
rect 22554 53564 22560 53576
rect 22515 53536 22560 53564
rect 2225 53527 2283 53533
rect 22554 53524 22560 53536
rect 22612 53524 22618 53576
rect 22738 53564 22744 53576
rect 22699 53536 22744 53564
rect 22738 53524 22744 53536
rect 22796 53524 22802 53576
rect 26786 53524 26792 53576
rect 26844 53564 26850 53576
rect 27249 53567 27307 53573
rect 27249 53564 27261 53567
rect 26844 53536 27261 53564
rect 26844 53524 26850 53536
rect 27249 53533 27261 53536
rect 27295 53533 27307 53567
rect 27249 53527 27307 53533
rect 27430 53524 27436 53576
rect 27488 53564 27494 53576
rect 28583 53567 28641 53573
rect 28583 53564 28595 53567
rect 27488 53536 28595 53564
rect 27488 53524 27494 53536
rect 28583 53533 28595 53536
rect 28629 53533 28641 53567
rect 28718 53564 28724 53576
rect 28679 53536 28724 53564
rect 28583 53527 28641 53533
rect 28718 53524 28724 53536
rect 28776 53524 28782 53576
rect 28813 53567 28871 53573
rect 28813 53533 28825 53567
rect 28859 53533 28871 53567
rect 28994 53564 29000 53576
rect 28955 53536 29000 53564
rect 28813 53527 28871 53533
rect 25406 53505 25412 53508
rect 25400 53459 25412 53505
rect 25464 53496 25470 53508
rect 25464 53468 25500 53496
rect 25406 53456 25412 53459
rect 25464 53456 25470 53468
rect 26878 53456 26884 53508
rect 26936 53496 26942 53508
rect 27341 53499 27399 53505
rect 27341 53496 27353 53499
rect 26936 53468 27353 53496
rect 26936 53456 26942 53468
rect 27341 53465 27353 53468
rect 27387 53465 27399 53499
rect 27341 53459 27399 53465
rect 28442 53456 28448 53508
rect 28500 53496 28506 53508
rect 28828 53496 28856 53527
rect 28994 53524 29000 53536
rect 29052 53524 29058 53576
rect 29546 53564 29552 53576
rect 29507 53536 29552 53564
rect 29546 53524 29552 53536
rect 29604 53524 29610 53576
rect 29638 53524 29644 53576
rect 29696 53564 29702 53576
rect 29805 53567 29863 53573
rect 29805 53564 29817 53567
rect 29696 53536 29817 53564
rect 29696 53524 29702 53536
rect 29805 53533 29817 53536
rect 29851 53533 29863 53567
rect 56318 53564 56324 53576
rect 56279 53536 56324 53564
rect 29805 53527 29863 53533
rect 56318 53524 56324 53536
rect 56376 53524 56382 53576
rect 28500 53468 30972 53496
rect 28500 53456 28506 53468
rect 22370 53388 22376 53440
rect 22428 53428 22434 53440
rect 22925 53431 22983 53437
rect 22925 53428 22937 53431
rect 22428 53400 22937 53428
rect 22428 53388 22434 53400
rect 22925 53397 22937 53400
rect 22971 53397 22983 53431
rect 22925 53391 22983 53397
rect 26513 53431 26571 53437
rect 26513 53397 26525 53431
rect 26559 53428 26571 53431
rect 27154 53428 27160 53440
rect 26559 53400 27160 53428
rect 26559 53397 26571 53400
rect 26513 53391 26571 53397
rect 27154 53388 27160 53400
rect 27212 53388 27218 53440
rect 30944 53437 30972 53468
rect 30929 53431 30987 53437
rect 30929 53397 30941 53431
rect 30975 53397 30987 53431
rect 30929 53391 30987 53397
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 25406 53224 25412 53236
rect 25367 53196 25412 53224
rect 25406 53184 25412 53196
rect 25464 53184 25470 53236
rect 27430 53224 27436 53236
rect 25516 53196 27200 53224
rect 27391 53196 27436 53224
rect 5166 53116 5172 53168
rect 5224 53156 5230 53168
rect 25516 53156 25544 53196
rect 5224 53128 25544 53156
rect 5224 53116 5230 53128
rect 25774 53116 25780 53168
rect 25832 53156 25838 53168
rect 27172 53156 27200 53196
rect 27430 53184 27436 53196
rect 27488 53184 27494 53236
rect 28166 53156 28172 53168
rect 25832 53128 26280 53156
rect 27172 53128 28172 53156
rect 25832 53116 25838 53128
rect 1946 53088 1952 53100
rect 1907 53060 1952 53088
rect 1946 53048 1952 53060
rect 2004 53048 2010 53100
rect 21821 53091 21879 53097
rect 21821 53057 21833 53091
rect 21867 53088 21879 53091
rect 21910 53088 21916 53100
rect 21867 53060 21916 53088
rect 21867 53057 21879 53060
rect 21821 53051 21879 53057
rect 21910 53048 21916 53060
rect 21968 53048 21974 53100
rect 22094 53097 22100 53100
rect 22088 53051 22100 53097
rect 22152 53088 22158 53100
rect 23658 53088 23664 53100
rect 22152 53060 22188 53088
rect 23619 53060 23664 53088
rect 22094 53048 22100 53051
rect 22152 53048 22158 53060
rect 23658 53048 23664 53060
rect 23716 53048 23722 53100
rect 23845 53091 23903 53097
rect 23845 53057 23857 53091
rect 23891 53088 23903 53091
rect 25498 53088 25504 53100
rect 23891 53060 25504 53088
rect 23891 53057 23903 53060
rect 23845 53051 23903 53057
rect 25498 53048 25504 53060
rect 25556 53048 25562 53100
rect 25593 53091 25651 53097
rect 25593 53057 25605 53091
rect 25639 53088 25651 53091
rect 26142 53088 26148 53100
rect 25639 53060 26148 53088
rect 25639 53057 25651 53060
rect 25593 53051 25651 53057
rect 26142 53048 26148 53060
rect 26200 53048 26206 53100
rect 26252 53097 26280 53128
rect 28166 53116 28172 53128
rect 28224 53116 28230 53168
rect 26237 53091 26295 53097
rect 26237 53057 26249 53091
rect 26283 53057 26295 53091
rect 26237 53051 26295 53057
rect 26878 53048 26884 53100
rect 26936 53088 26942 53100
rect 26973 53091 27031 53097
rect 26973 53088 26985 53091
rect 26936 53060 26985 53088
rect 26936 53048 26942 53060
rect 26973 53057 26985 53060
rect 27019 53057 27031 53091
rect 27246 53088 27252 53100
rect 27207 53060 27252 53088
rect 26973 53051 27031 53057
rect 27246 53048 27252 53060
rect 27304 53048 27310 53100
rect 27338 53048 27344 53100
rect 27396 53088 27402 53100
rect 28077 53091 28135 53097
rect 28077 53088 28089 53091
rect 27396 53060 28089 53088
rect 27396 53048 27402 53060
rect 28077 53057 28089 53060
rect 28123 53057 28135 53091
rect 28077 53051 28135 53057
rect 56318 53048 56324 53100
rect 56376 53088 56382 53100
rect 58069 53091 58127 53097
rect 58069 53088 58081 53091
rect 56376 53060 58081 53088
rect 56376 53048 56382 53060
rect 58069 53057 58081 53060
rect 58115 53057 58127 53091
rect 58069 53051 58127 53057
rect 2133 53023 2191 53029
rect 2133 52989 2145 53023
rect 2179 53020 2191 53023
rect 2406 53020 2412 53032
rect 2179 52992 2412 53020
rect 2179 52989 2191 52992
rect 2133 52983 2191 52989
rect 2406 52980 2412 52992
rect 2464 52980 2470 53032
rect 2774 53020 2780 53032
rect 2735 52992 2780 53020
rect 2774 52980 2780 52992
rect 2832 52980 2838 53032
rect 26053 53023 26111 53029
rect 26053 52989 26065 53023
rect 26099 53020 26111 53023
rect 26099 52992 26234 53020
rect 26099 52989 26111 52992
rect 26053 52983 26111 52989
rect 26206 52952 26234 52992
rect 26786 52980 26792 53032
rect 26844 53020 26850 53032
rect 27065 53023 27123 53029
rect 27065 53020 27077 53023
rect 26844 52992 27077 53020
rect 26844 52980 26850 52992
rect 27065 52989 27077 52992
rect 27111 52989 27123 53023
rect 27065 52983 27123 52989
rect 27154 52952 27160 52964
rect 26206 52924 27160 52952
rect 23198 52884 23204 52896
rect 23159 52856 23204 52884
rect 23198 52844 23204 52856
rect 23256 52844 23262 52896
rect 23474 52844 23480 52896
rect 23532 52884 23538 52896
rect 24029 52887 24087 52893
rect 24029 52884 24041 52887
rect 23532 52856 24041 52884
rect 23532 52844 23538 52856
rect 24029 52853 24041 52856
rect 24075 52853 24087 52887
rect 26418 52884 26424 52896
rect 26379 52856 26424 52884
rect 24029 52847 24087 52853
rect 26418 52844 26424 52856
rect 26476 52844 26482 52896
rect 26988 52893 27016 52924
rect 27154 52912 27160 52924
rect 27212 52912 27218 52964
rect 26973 52887 27031 52893
rect 26973 52853 26985 52887
rect 27019 52853 27031 52887
rect 26973 52847 27031 52853
rect 27062 52844 27068 52896
rect 27120 52884 27126 52896
rect 27893 52887 27951 52893
rect 27893 52884 27905 52887
rect 27120 52856 27905 52884
rect 27120 52844 27126 52856
rect 27893 52853 27905 52856
rect 27939 52853 27951 52887
rect 27893 52847 27951 52853
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 2406 52680 2412 52692
rect 2367 52652 2412 52680
rect 2406 52640 2412 52652
rect 2464 52640 2470 52692
rect 21453 52615 21511 52621
rect 21453 52581 21465 52615
rect 21499 52612 21511 52615
rect 22094 52612 22100 52624
rect 21499 52584 22100 52612
rect 21499 52581 21511 52584
rect 21453 52575 21511 52581
rect 22094 52572 22100 52584
rect 22152 52572 22158 52624
rect 26878 52612 26884 52624
rect 26839 52584 26884 52612
rect 26878 52572 26884 52584
rect 26936 52572 26942 52624
rect 25038 52504 25044 52556
rect 25096 52544 25102 52556
rect 25501 52547 25559 52553
rect 25501 52544 25513 52547
rect 25096 52516 25513 52544
rect 25096 52504 25102 52516
rect 25501 52513 25513 52516
rect 25547 52513 25559 52547
rect 25501 52507 25559 52513
rect 2314 52476 2320 52488
rect 2275 52448 2320 52476
rect 2314 52436 2320 52448
rect 2372 52436 2378 52488
rect 3142 52476 3148 52488
rect 3103 52448 3148 52476
rect 3142 52436 3148 52448
rect 3200 52436 3206 52488
rect 3789 52479 3847 52485
rect 3789 52445 3801 52479
rect 3835 52476 3847 52479
rect 5166 52476 5172 52488
rect 3835 52448 5172 52476
rect 3835 52445 3847 52448
rect 3789 52439 3847 52445
rect 5166 52436 5172 52448
rect 5224 52436 5230 52488
rect 21637 52479 21695 52485
rect 21637 52445 21649 52479
rect 21683 52476 21695 52479
rect 21683 52448 21864 52476
rect 21683 52445 21695 52448
rect 21637 52439 21695 52445
rect 21836 52408 21864 52448
rect 21910 52436 21916 52488
rect 21968 52476 21974 52488
rect 22097 52479 22155 52485
rect 22097 52476 22109 52479
rect 21968 52448 22109 52476
rect 21968 52436 21974 52448
rect 22097 52445 22109 52448
rect 22143 52476 22155 52479
rect 25056 52476 25084 52504
rect 22143 52448 25084 52476
rect 25768 52479 25826 52485
rect 22143 52445 22155 52448
rect 22097 52439 22155 52445
rect 25768 52445 25780 52479
rect 25814 52476 25826 52479
rect 26970 52476 26976 52488
rect 25814 52448 26976 52476
rect 25814 52445 25826 52448
rect 25768 52439 25826 52445
rect 26970 52436 26976 52448
rect 27028 52436 27034 52488
rect 28994 52436 29000 52488
rect 29052 52476 29058 52488
rect 30190 52476 30196 52488
rect 29052 52448 30196 52476
rect 29052 52436 29058 52448
rect 30190 52436 30196 52448
rect 30248 52436 30254 52488
rect 22364 52411 22422 52417
rect 21836 52380 22324 52408
rect 3878 52340 3884 52352
rect 3839 52312 3884 52340
rect 3878 52300 3884 52312
rect 3936 52300 3942 52352
rect 22296 52340 22324 52380
rect 22364 52377 22376 52411
rect 22410 52408 22422 52411
rect 22462 52408 22468 52420
rect 22410 52380 22468 52408
rect 22410 52377 22422 52380
rect 22364 52371 22422 52377
rect 22462 52368 22468 52380
rect 22520 52368 22526 52420
rect 22646 52340 22652 52352
rect 22296 52312 22652 52340
rect 22646 52300 22652 52312
rect 22704 52300 22710 52352
rect 23477 52343 23535 52349
rect 23477 52309 23489 52343
rect 23523 52340 23535 52343
rect 23750 52340 23756 52352
rect 23523 52312 23756 52340
rect 23523 52309 23535 52312
rect 23477 52303 23535 52309
rect 23750 52300 23756 52312
rect 23808 52300 23814 52352
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 22554 52096 22560 52148
rect 22612 52136 22618 52148
rect 23106 52136 23112 52148
rect 22612 52108 23112 52136
rect 22612 52096 22618 52108
rect 23106 52096 23112 52108
rect 23164 52136 23170 52148
rect 23293 52139 23351 52145
rect 23293 52136 23305 52139
rect 23164 52108 23305 52136
rect 23164 52096 23170 52108
rect 23293 52105 23305 52108
rect 23339 52105 23351 52139
rect 23293 52099 23351 52105
rect 2409 52071 2467 52077
rect 2409 52037 2421 52071
rect 2455 52068 2467 52071
rect 3878 52068 3884 52080
rect 2455 52040 3884 52068
rect 2455 52037 2467 52040
rect 2409 52031 2467 52037
rect 3878 52028 3884 52040
rect 3936 52028 3942 52080
rect 20257 52071 20315 52077
rect 20257 52068 20269 52071
rect 19444 52040 20269 52068
rect 19444 52009 19472 52040
rect 20257 52037 20269 52040
rect 20303 52037 20315 52071
rect 20257 52031 20315 52037
rect 22094 52028 22100 52080
rect 22152 52077 22158 52080
rect 22152 52071 22216 52077
rect 22152 52037 22170 52071
rect 22204 52037 22216 52071
rect 23308 52068 23336 52099
rect 23658 52096 23664 52148
rect 23716 52136 23722 52148
rect 23937 52139 23995 52145
rect 23937 52136 23949 52139
rect 23716 52108 23949 52136
rect 23716 52096 23722 52108
rect 23937 52105 23949 52108
rect 23983 52105 23995 52139
rect 23937 52099 23995 52105
rect 26421 52139 26479 52145
rect 26421 52105 26433 52139
rect 26467 52136 26479 52139
rect 26786 52136 26792 52148
rect 26467 52108 26792 52136
rect 26467 52105 26479 52108
rect 26421 52099 26479 52105
rect 26786 52096 26792 52108
rect 26844 52096 26850 52148
rect 26970 52136 26976 52148
rect 26931 52108 26976 52136
rect 26970 52096 26976 52108
rect 27028 52096 27034 52148
rect 24121 52071 24179 52077
rect 24121 52068 24133 52071
rect 23308 52040 24133 52068
rect 22152 52031 22216 52037
rect 24121 52037 24133 52040
rect 24167 52037 24179 52071
rect 24121 52031 24179 52037
rect 25308 52071 25366 52077
rect 25308 52037 25320 52071
rect 25354 52068 25366 52071
rect 27062 52068 27068 52080
rect 25354 52040 27068 52068
rect 25354 52037 25366 52040
rect 25308 52031 25366 52037
rect 22152 52028 22158 52031
rect 27062 52028 27068 52040
rect 27120 52028 27126 52080
rect 32122 52068 32128 52080
rect 30208 52040 32128 52068
rect 19429 52003 19487 52009
rect 19429 51969 19441 52003
rect 19475 51969 19487 52003
rect 19978 52000 19984 52012
rect 19939 51972 19984 52000
rect 19429 51963 19487 51969
rect 19978 51960 19984 51972
rect 20036 51960 20042 52012
rect 20070 51960 20076 52012
rect 20128 52000 20134 52012
rect 21910 52000 21916 52012
rect 20128 51972 20173 52000
rect 21871 51972 21916 52000
rect 20128 51960 20134 51972
rect 21910 51960 21916 51972
rect 21968 51960 21974 52012
rect 23198 51960 23204 52012
rect 23256 52000 23262 52012
rect 24029 52003 24087 52009
rect 24029 52000 24041 52003
rect 23256 51972 24041 52000
rect 23256 51960 23262 51972
rect 24029 51969 24041 51972
rect 24075 51969 24087 52003
rect 25038 52000 25044 52012
rect 24999 51972 25044 52000
rect 24029 51963 24087 51969
rect 25038 51960 25044 51972
rect 25096 51960 25102 52012
rect 26418 51960 26424 52012
rect 26476 52000 26482 52012
rect 27157 52003 27215 52009
rect 27157 52000 27169 52003
rect 26476 51972 27169 52000
rect 26476 51960 26482 51972
rect 27157 51969 27169 51972
rect 27203 51969 27215 52003
rect 27157 51963 27215 51969
rect 28994 51960 29000 52012
rect 29052 52000 29058 52012
rect 29546 52000 29552 52012
rect 29052 51972 29552 52000
rect 29052 51960 29058 51972
rect 29546 51960 29552 51972
rect 29604 52000 29610 52012
rect 30208 52009 30236 52040
rect 32122 52028 32128 52040
rect 32180 52028 32186 52080
rect 30466 52009 30472 52012
rect 30193 52003 30251 52009
rect 30193 52000 30205 52003
rect 29604 51972 30205 52000
rect 29604 51960 29610 51972
rect 30193 51969 30205 51972
rect 30239 51969 30251 52003
rect 30193 51963 30251 51969
rect 30460 51963 30472 52009
rect 30524 52000 30530 52012
rect 30524 51972 30560 52000
rect 30466 51960 30472 51963
rect 30524 51960 30530 51972
rect 31386 51960 31392 52012
rect 31444 52000 31450 52012
rect 32309 52003 32367 52009
rect 32309 52000 32321 52003
rect 31444 51972 32321 52000
rect 31444 51960 31450 51972
rect 32309 51969 32321 51972
rect 32355 51969 32367 52003
rect 32309 51963 32367 51969
rect 32493 52003 32551 52009
rect 32493 51969 32505 52003
rect 32539 52000 32551 52003
rect 33137 52003 33195 52009
rect 33137 52000 33149 52003
rect 32539 51972 33149 52000
rect 32539 51969 32551 51972
rect 32493 51963 32551 51969
rect 33137 51969 33149 51972
rect 33183 51969 33195 52003
rect 33137 51963 33195 51969
rect 2225 51935 2283 51941
rect 2225 51901 2237 51935
rect 2271 51932 2283 51935
rect 3142 51932 3148 51944
rect 2271 51904 3148 51932
rect 2271 51901 2283 51904
rect 2225 51895 2283 51901
rect 3142 51892 3148 51904
rect 3200 51892 3206 51944
rect 3234 51892 3240 51944
rect 3292 51932 3298 51944
rect 32125 51935 32183 51941
rect 3292 51904 3337 51932
rect 3292 51892 3298 51904
rect 32125 51901 32137 51935
rect 32171 51932 32183 51935
rect 32398 51932 32404 51944
rect 32171 51904 32404 51932
rect 32171 51901 32183 51904
rect 32125 51895 32183 51901
rect 23750 51864 23756 51876
rect 23711 51836 23756 51864
rect 23750 51824 23756 51836
rect 23808 51824 23814 51876
rect 31573 51867 31631 51873
rect 31573 51833 31585 51867
rect 31619 51864 31631 51867
rect 32140 51864 32168 51895
rect 32398 51892 32404 51904
rect 32456 51892 32462 51944
rect 31619 51836 32168 51864
rect 31619 51833 31631 51836
rect 31573 51827 31631 51833
rect 19245 51799 19303 51805
rect 19245 51765 19257 51799
rect 19291 51796 19303 51799
rect 19334 51796 19340 51808
rect 19291 51768 19340 51796
rect 19291 51765 19303 51768
rect 19245 51759 19303 51765
rect 19334 51756 19340 51768
rect 19392 51756 19398 51808
rect 24210 51756 24216 51808
rect 24268 51796 24274 51808
rect 24305 51799 24363 51805
rect 24305 51796 24317 51799
rect 24268 51768 24317 51796
rect 24268 51756 24274 51768
rect 24305 51765 24317 51768
rect 24351 51765 24363 51799
rect 24305 51759 24363 51765
rect 32306 51756 32312 51808
rect 32364 51796 32370 51808
rect 32953 51799 33011 51805
rect 32953 51796 32965 51799
rect 32364 51768 32965 51796
rect 32364 51756 32370 51768
rect 32953 51765 32965 51768
rect 32999 51765 33011 51799
rect 32953 51759 33011 51765
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 21637 51595 21695 51601
rect 21637 51561 21649 51595
rect 21683 51592 21695 51595
rect 22186 51592 22192 51604
rect 21683 51564 22192 51592
rect 21683 51561 21695 51564
rect 21637 51555 21695 51561
rect 22186 51552 22192 51564
rect 22244 51552 22250 51604
rect 22646 51592 22652 51604
rect 22607 51564 22652 51592
rect 22646 51552 22652 51564
rect 22704 51552 22710 51604
rect 23385 51595 23443 51601
rect 23385 51561 23397 51595
rect 23431 51592 23443 51595
rect 23658 51592 23664 51604
rect 23431 51564 23664 51592
rect 23431 51561 23443 51564
rect 23385 51555 23443 51561
rect 23658 51552 23664 51564
rect 23716 51552 23722 51604
rect 25961 51595 26019 51601
rect 25961 51561 25973 51595
rect 26007 51592 26019 51595
rect 27338 51592 27344 51604
rect 26007 51564 27344 51592
rect 26007 51561 26019 51564
rect 25961 51555 26019 51561
rect 27338 51552 27344 51564
rect 27396 51552 27402 51604
rect 30466 51552 30472 51604
rect 30524 51592 30530 51604
rect 30561 51595 30619 51601
rect 30561 51592 30573 51595
rect 30524 51564 30573 51592
rect 30524 51552 30530 51564
rect 30561 51561 30573 51564
rect 30607 51561 30619 51595
rect 30561 51555 30619 51561
rect 22281 51459 22339 51465
rect 22281 51425 22293 51459
rect 22327 51456 22339 51459
rect 22327 51428 23152 51456
rect 22327 51425 22339 51428
rect 22281 51419 22339 51425
rect 19242 51388 19248 51400
rect 19203 51360 19248 51388
rect 19242 51348 19248 51360
rect 19300 51348 19306 51400
rect 19334 51348 19340 51400
rect 19392 51388 19398 51400
rect 19501 51391 19559 51397
rect 19501 51388 19513 51391
rect 19392 51360 19513 51388
rect 19392 51348 19398 51360
rect 19501 51357 19513 51360
rect 19547 51357 19559 51391
rect 19501 51351 19559 51357
rect 21821 51391 21879 51397
rect 21821 51357 21833 51391
rect 21867 51388 21879 51391
rect 22370 51388 22376 51400
rect 21867 51360 22376 51388
rect 21867 51357 21879 51360
rect 21821 51351 21879 51357
rect 22370 51348 22376 51360
rect 22428 51348 22434 51400
rect 22465 51391 22523 51397
rect 22465 51357 22477 51391
rect 22511 51388 22523 51391
rect 22738 51388 22744 51400
rect 22511 51360 22744 51388
rect 22511 51357 22523 51360
rect 22465 51351 22523 51357
rect 22738 51348 22744 51360
rect 22796 51348 22802 51400
rect 23124 51388 23152 51428
rect 23198 51416 23204 51468
rect 23256 51456 23262 51468
rect 25593 51459 25651 51465
rect 23256 51428 23301 51456
rect 23256 51416 23262 51428
rect 25593 51425 25605 51459
rect 25639 51456 25651 51459
rect 26878 51456 26884 51468
rect 25639 51428 26884 51456
rect 25639 51425 25651 51428
rect 25593 51419 25651 51425
rect 26878 51416 26884 51428
rect 26936 51416 26942 51468
rect 29932 51428 31432 51456
rect 23385 51391 23443 51397
rect 23385 51388 23397 51391
rect 23124 51360 23397 51388
rect 23385 51357 23397 51360
rect 23431 51388 23443 51391
rect 23750 51388 23756 51400
rect 23431 51360 23756 51388
rect 23431 51357 23443 51360
rect 23385 51351 23443 51357
rect 23750 51348 23756 51360
rect 23808 51348 23814 51400
rect 25774 51388 25780 51400
rect 25735 51360 25780 51388
rect 25774 51348 25780 51360
rect 25832 51348 25838 51400
rect 28997 51391 29055 51397
rect 28997 51357 29009 51391
rect 29043 51388 29055 51391
rect 29638 51388 29644 51400
rect 29043 51360 29644 51388
rect 29043 51357 29055 51360
rect 28997 51351 29055 51357
rect 29638 51348 29644 51360
rect 29696 51348 29702 51400
rect 29730 51348 29736 51400
rect 29788 51388 29794 51400
rect 29932 51397 29960 51428
rect 31404 51400 31432 51428
rect 29917 51391 29975 51397
rect 29788 51360 29833 51388
rect 29788 51348 29794 51360
rect 29917 51357 29929 51391
rect 29963 51357 29975 51391
rect 29917 51351 29975 51357
rect 30101 51391 30159 51397
rect 30101 51357 30113 51391
rect 30147 51388 30159 51391
rect 30745 51391 30803 51397
rect 30745 51388 30757 51391
rect 30147 51360 30757 51388
rect 30147 51357 30159 51360
rect 30101 51351 30159 51357
rect 30745 51357 30757 51360
rect 30791 51357 30803 51391
rect 30745 51351 30803 51357
rect 31297 51391 31355 51397
rect 31297 51357 31309 51391
rect 31343 51357 31355 51391
rect 31297 51351 31355 51357
rect 23106 51320 23112 51332
rect 23067 51292 23112 51320
rect 23106 51280 23112 51292
rect 23164 51280 23170 51332
rect 25498 51280 25504 51332
rect 25556 51320 25562 51332
rect 29932 51320 29960 51351
rect 25556 51292 29960 51320
rect 31312 51320 31340 51351
rect 31386 51348 31392 51400
rect 31444 51388 31450 51400
rect 32033 51391 32091 51397
rect 31444 51360 31537 51388
rect 31444 51348 31450 51360
rect 32033 51357 32045 51391
rect 32079 51388 32091 51391
rect 32122 51388 32128 51400
rect 32079 51360 32128 51388
rect 32079 51357 32091 51360
rect 32033 51351 32091 51357
rect 32122 51348 32128 51360
rect 32180 51348 32186 51400
rect 32306 51397 32312 51400
rect 32300 51388 32312 51397
rect 32267 51360 32312 51388
rect 32300 51351 32312 51360
rect 32306 51348 32312 51351
rect 32364 51348 32370 51400
rect 32582 51348 32588 51400
rect 32640 51388 32646 51400
rect 34057 51391 34115 51397
rect 34057 51388 34069 51391
rect 32640 51360 34069 51388
rect 32640 51348 32646 51360
rect 34057 51357 34069 51360
rect 34103 51357 34115 51391
rect 34057 51351 34115 51357
rect 36170 51348 36176 51400
rect 36228 51388 36234 51400
rect 56965 51391 57023 51397
rect 56965 51388 56977 51391
rect 36228 51360 56977 51388
rect 36228 51348 36234 51360
rect 56965 51357 56977 51360
rect 57011 51388 57023 51391
rect 57514 51388 57520 51400
rect 57011 51360 57520 51388
rect 57011 51357 57023 51360
rect 56965 51351 57023 51357
rect 57514 51348 57520 51360
rect 57572 51348 57578 51400
rect 57790 51388 57796 51400
rect 57751 51360 57796 51388
rect 57790 51348 57796 51360
rect 57848 51348 57854 51400
rect 32490 51320 32496 51332
rect 31312 51292 32496 51320
rect 25556 51280 25562 51292
rect 32490 51280 32496 51292
rect 32548 51320 32554 51332
rect 33134 51320 33140 51332
rect 32548 51292 33140 51320
rect 32548 51280 32554 51292
rect 33134 51280 33140 51292
rect 33192 51280 33198 51332
rect 20622 51252 20628 51264
rect 20583 51224 20628 51252
rect 20622 51212 20628 51224
rect 20680 51212 20686 51264
rect 23569 51255 23627 51261
rect 23569 51221 23581 51255
rect 23615 51252 23627 51255
rect 24578 51252 24584 51264
rect 23615 51224 24584 51252
rect 23615 51221 23627 51224
rect 23569 51215 23627 51221
rect 24578 51212 24584 51224
rect 24636 51212 24642 51264
rect 28810 51252 28816 51264
rect 28771 51224 28816 51252
rect 28810 51212 28816 51224
rect 28868 51212 28874 51264
rect 31573 51255 31631 51261
rect 31573 51221 31585 51255
rect 31619 51252 31631 51255
rect 33042 51252 33048 51264
rect 31619 51224 33048 51252
rect 31619 51221 31631 51224
rect 31573 51215 31631 51221
rect 33042 51212 33048 51224
rect 33100 51212 33106 51264
rect 33410 51252 33416 51264
rect 33371 51224 33416 51252
rect 33410 51212 33416 51224
rect 33468 51212 33474 51264
rect 33870 51252 33876 51264
rect 33831 51224 33876 51252
rect 33870 51212 33876 51224
rect 33928 51212 33934 51264
rect 57054 51252 57060 51264
rect 57015 51224 57060 51252
rect 57054 51212 57060 51224
rect 57112 51212 57118 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 22462 51008 22468 51060
rect 22520 51048 22526 51060
rect 23293 51051 23351 51057
rect 23293 51048 23305 51051
rect 22520 51020 23305 51048
rect 22520 51008 22526 51020
rect 23293 51017 23305 51020
rect 23339 51017 23351 51051
rect 23293 51011 23351 51017
rect 31573 51051 31631 51057
rect 31573 51017 31585 51051
rect 31619 51048 31631 51051
rect 32582 51048 32588 51060
rect 31619 51020 32588 51048
rect 31619 51017 31631 51020
rect 31573 51011 31631 51017
rect 32582 51008 32588 51020
rect 32640 51008 32646 51060
rect 33134 51008 33140 51060
rect 33192 51048 33198 51060
rect 33505 51051 33563 51057
rect 33505 51048 33517 51051
rect 33192 51020 33517 51048
rect 33192 51008 33198 51020
rect 33505 51017 33517 51020
rect 33551 51048 33563 51051
rect 33551 51020 34008 51048
rect 33551 51017 33563 51020
rect 33505 51011 33563 51017
rect 20254 50980 20260 50992
rect 19812 50952 20260 50980
rect 19812 50921 19840 50952
rect 20254 50940 20260 50952
rect 20312 50980 20318 50992
rect 20622 50980 20628 50992
rect 20312 50952 20628 50980
rect 20312 50940 20318 50952
rect 20622 50940 20628 50952
rect 20680 50940 20686 50992
rect 23198 50980 23204 50992
rect 22572 50952 23204 50980
rect 19797 50915 19855 50921
rect 19797 50881 19809 50915
rect 19843 50881 19855 50915
rect 19797 50875 19855 50881
rect 19889 50915 19947 50921
rect 19889 50881 19901 50915
rect 19935 50912 19947 50915
rect 20070 50912 20076 50924
rect 19935 50884 20076 50912
rect 19935 50881 19947 50884
rect 19889 50875 19947 50881
rect 20070 50872 20076 50884
rect 20128 50912 20134 50924
rect 22572 50921 22600 50952
rect 23198 50940 23204 50952
rect 23256 50940 23262 50992
rect 28902 50980 28908 50992
rect 28552 50952 28908 50980
rect 22557 50915 22615 50921
rect 20128 50884 22094 50912
rect 20128 50872 20134 50884
rect 22066 50776 22094 50884
rect 22557 50881 22569 50915
rect 22603 50881 22615 50915
rect 22557 50875 22615 50881
rect 22649 50915 22707 50921
rect 22649 50881 22661 50915
rect 22695 50881 22707 50915
rect 23474 50912 23480 50924
rect 23435 50884 23480 50912
rect 22649 50875 22707 50881
rect 22664 50844 22692 50875
rect 23474 50872 23480 50884
rect 23532 50872 23538 50924
rect 24949 50915 25007 50921
rect 24949 50881 24961 50915
rect 24995 50881 25007 50915
rect 24949 50875 25007 50881
rect 22738 50844 22744 50856
rect 22651 50816 22744 50844
rect 22738 50804 22744 50816
rect 22796 50844 22802 50856
rect 24964 50844 24992 50875
rect 25498 50872 25504 50924
rect 25556 50912 25562 50924
rect 25685 50915 25743 50921
rect 25685 50912 25697 50915
rect 25556 50884 25697 50912
rect 25556 50872 25562 50884
rect 25685 50881 25697 50884
rect 25731 50881 25743 50915
rect 25685 50875 25743 50881
rect 28258 50872 28264 50924
rect 28316 50912 28322 50924
rect 28552 50921 28580 50952
rect 28902 50940 28908 50952
rect 28960 50940 28966 50992
rect 29454 50940 29460 50992
rect 29512 50980 29518 50992
rect 30377 50983 30435 50989
rect 30377 50980 30389 50983
rect 29512 50952 30389 50980
rect 29512 50940 29518 50952
rect 30377 50949 30389 50952
rect 30423 50949 30435 50983
rect 30377 50943 30435 50949
rect 30593 50983 30651 50989
rect 30593 50949 30605 50983
rect 30639 50980 30651 50983
rect 32392 50983 32450 50989
rect 30639 50952 31754 50980
rect 30639 50949 30651 50952
rect 30593 50943 30651 50949
rect 28810 50921 28816 50924
rect 28537 50915 28595 50921
rect 28537 50912 28549 50915
rect 28316 50884 28549 50912
rect 28316 50872 28322 50884
rect 28537 50881 28549 50884
rect 28583 50881 28595 50915
rect 28804 50912 28816 50921
rect 28771 50884 28816 50912
rect 28537 50875 28595 50881
rect 28804 50875 28816 50884
rect 28810 50872 28816 50875
rect 28868 50872 28874 50924
rect 31386 50912 31392 50924
rect 31347 50884 31392 50912
rect 31386 50872 31392 50884
rect 31444 50872 31450 50924
rect 31726 50912 31754 50952
rect 32392 50949 32404 50983
rect 32438 50980 32450 50983
rect 33870 50980 33876 50992
rect 32438 50952 33876 50980
rect 32438 50949 32450 50952
rect 32392 50943 32450 50949
rect 33870 50940 33876 50952
rect 33928 50940 33934 50992
rect 33980 50989 34008 51020
rect 33965 50983 34023 50989
rect 33965 50949 33977 50983
rect 34011 50949 34023 50983
rect 33965 50943 34023 50949
rect 32674 50912 32680 50924
rect 31726 50884 32680 50912
rect 32674 50872 32680 50884
rect 32732 50872 32738 50924
rect 33318 50872 33324 50924
rect 33376 50912 33382 50924
rect 34241 50915 34299 50921
rect 34241 50912 34253 50915
rect 33376 50884 34253 50912
rect 33376 50872 33382 50884
rect 34241 50881 34253 50884
rect 34287 50881 34299 50915
rect 34241 50875 34299 50881
rect 25409 50847 25467 50853
rect 25409 50844 25421 50847
rect 22796 50816 24808 50844
rect 24964 50816 25421 50844
rect 22796 50804 22802 50816
rect 23492 50788 23520 50816
rect 22066 50748 23428 50776
rect 18690 50668 18696 50720
rect 18748 50708 18754 50720
rect 20073 50711 20131 50717
rect 20073 50708 20085 50711
rect 18748 50680 20085 50708
rect 18748 50668 18754 50680
rect 20073 50677 20085 50680
rect 20119 50677 20131 50711
rect 20073 50671 20131 50677
rect 22370 50668 22376 50720
rect 22428 50708 22434 50720
rect 22833 50711 22891 50717
rect 22833 50708 22845 50711
rect 22428 50680 22845 50708
rect 22428 50668 22434 50680
rect 22833 50677 22845 50680
rect 22879 50677 22891 50711
rect 23400 50708 23428 50748
rect 23474 50736 23480 50788
rect 23532 50736 23538 50788
rect 24780 50785 24808 50816
rect 25409 50813 25421 50816
rect 25455 50844 25467 50847
rect 25590 50844 25596 50856
rect 25455 50816 25596 50844
rect 25455 50813 25467 50816
rect 25409 50807 25467 50813
rect 25590 50804 25596 50816
rect 25648 50804 25654 50856
rect 31205 50847 31263 50853
rect 31205 50813 31217 50847
rect 31251 50844 31263 50847
rect 31662 50844 31668 50856
rect 31251 50816 31668 50844
rect 31251 50813 31263 50816
rect 31205 50807 31263 50813
rect 31662 50804 31668 50816
rect 31720 50844 31726 50856
rect 31938 50844 31944 50856
rect 31720 50816 31944 50844
rect 31720 50804 31726 50816
rect 31938 50804 31944 50816
rect 31996 50804 32002 50856
rect 32122 50844 32128 50856
rect 32083 50816 32128 50844
rect 32122 50804 32128 50816
rect 32180 50804 32186 50856
rect 33502 50804 33508 50856
rect 33560 50844 33566 50856
rect 34057 50847 34115 50853
rect 34057 50844 34069 50847
rect 33560 50816 34069 50844
rect 33560 50804 33566 50816
rect 34057 50813 34069 50816
rect 34103 50813 34115 50847
rect 34057 50807 34115 50813
rect 24765 50779 24823 50785
rect 24765 50745 24777 50779
rect 24811 50745 24823 50779
rect 24765 50739 24823 50745
rect 29822 50736 29828 50788
rect 29880 50776 29886 50788
rect 34425 50779 34483 50785
rect 34425 50776 34437 50779
rect 29880 50748 31754 50776
rect 29880 50736 29886 50748
rect 25774 50708 25780 50720
rect 23400 50680 25780 50708
rect 22833 50671 22891 50677
rect 25774 50668 25780 50680
rect 25832 50668 25838 50720
rect 29730 50668 29736 50720
rect 29788 50708 29794 50720
rect 29917 50711 29975 50717
rect 29917 50708 29929 50711
rect 29788 50680 29929 50708
rect 29788 50668 29794 50680
rect 29917 50677 29929 50680
rect 29963 50708 29975 50711
rect 30561 50711 30619 50717
rect 30561 50708 30573 50711
rect 29963 50680 30573 50708
rect 29963 50677 29975 50680
rect 29917 50671 29975 50677
rect 30561 50677 30573 50680
rect 30607 50677 30619 50711
rect 30561 50671 30619 50677
rect 30745 50711 30803 50717
rect 30745 50677 30757 50711
rect 30791 50708 30803 50711
rect 30834 50708 30840 50720
rect 30791 50680 30840 50708
rect 30791 50677 30803 50680
rect 30745 50671 30803 50677
rect 30834 50668 30840 50680
rect 30892 50668 30898 50720
rect 31726 50708 31754 50748
rect 33060 50748 34437 50776
rect 33060 50708 33088 50748
rect 34425 50745 34437 50748
rect 34471 50745 34483 50779
rect 34425 50739 34483 50745
rect 33962 50708 33968 50720
rect 31726 50680 33088 50708
rect 33923 50680 33968 50708
rect 33962 50668 33968 50680
rect 34020 50668 34026 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 25038 50504 25044 50516
rect 24999 50476 25044 50504
rect 25038 50464 25044 50476
rect 25096 50464 25102 50516
rect 30653 50507 30711 50513
rect 30653 50504 30665 50507
rect 28920 50476 30665 50504
rect 19242 50368 19248 50380
rect 19203 50340 19248 50368
rect 19242 50328 19248 50340
rect 19300 50328 19306 50380
rect 26050 50328 26056 50380
rect 26108 50368 26114 50380
rect 26145 50371 26203 50377
rect 26145 50368 26157 50371
rect 26108 50340 26157 50368
rect 26108 50328 26114 50340
rect 26145 50337 26157 50340
rect 26191 50337 26203 50371
rect 26145 50331 26203 50337
rect 18690 50300 18696 50312
rect 18651 50272 18696 50300
rect 18690 50260 18696 50272
rect 18748 50260 18754 50312
rect 22370 50300 22376 50312
rect 22331 50272 22376 50300
rect 22370 50260 22376 50272
rect 22428 50260 22434 50312
rect 25590 50260 25596 50312
rect 25648 50300 25654 50312
rect 25869 50303 25927 50309
rect 25869 50300 25881 50303
rect 25648 50272 25881 50300
rect 25648 50260 25654 50272
rect 25869 50269 25881 50272
rect 25915 50269 25927 50303
rect 25869 50263 25927 50269
rect 27617 50303 27675 50309
rect 27617 50269 27629 50303
rect 27663 50300 27675 50303
rect 28258 50300 28264 50312
rect 27663 50272 28264 50300
rect 27663 50269 27675 50272
rect 27617 50263 27675 50269
rect 28258 50260 28264 50272
rect 28316 50260 28322 50312
rect 19490 50235 19548 50241
rect 19490 50232 19502 50235
rect 18524 50204 19502 50232
rect 18524 50173 18552 50204
rect 19490 50201 19502 50204
rect 19536 50201 19548 50235
rect 19490 50195 19548 50201
rect 24949 50235 25007 50241
rect 24949 50201 24961 50235
rect 24995 50232 25007 50235
rect 25958 50232 25964 50244
rect 24995 50204 25964 50232
rect 24995 50201 25007 50204
rect 24949 50195 25007 50201
rect 25958 50192 25964 50204
rect 26016 50192 26022 50244
rect 27884 50235 27942 50241
rect 27884 50201 27896 50235
rect 27930 50232 27942 50235
rect 28920 50232 28948 50476
rect 30653 50473 30665 50476
rect 30699 50473 30711 50507
rect 30653 50467 30711 50473
rect 31938 50464 31944 50516
rect 31996 50504 32002 50516
rect 33318 50504 33324 50516
rect 31996 50476 33324 50504
rect 31996 50464 32002 50476
rect 33318 50464 33324 50476
rect 33376 50464 33382 50516
rect 33502 50504 33508 50516
rect 33463 50476 33508 50504
rect 33502 50464 33508 50476
rect 33560 50464 33566 50516
rect 28997 50439 29055 50445
rect 28997 50405 29009 50439
rect 29043 50405 29055 50439
rect 28997 50399 29055 50405
rect 29549 50439 29607 50445
rect 29549 50405 29561 50439
rect 29595 50436 29607 50439
rect 57790 50436 57796 50448
rect 29595 50408 31156 50436
rect 29595 50405 29607 50408
rect 29549 50399 29607 50405
rect 29012 50368 29040 50399
rect 30834 50368 30840 50380
rect 29012 50340 30052 50368
rect 30795 50340 30840 50368
rect 30024 50312 30052 50340
rect 30834 50328 30840 50340
rect 30892 50328 30898 50380
rect 31128 50377 31156 50408
rect 56336 50408 57796 50436
rect 56336 50377 56364 50408
rect 57790 50396 57796 50408
rect 57848 50396 57854 50448
rect 31113 50371 31171 50377
rect 31113 50337 31125 50371
rect 31159 50337 31171 50371
rect 31113 50331 31171 50337
rect 56321 50371 56379 50377
rect 56321 50337 56333 50371
rect 56367 50337 56379 50371
rect 56321 50331 56379 50337
rect 56505 50371 56563 50377
rect 56505 50337 56517 50371
rect 56551 50368 56563 50371
rect 57054 50368 57060 50380
rect 56551 50340 57060 50368
rect 56551 50337 56563 50340
rect 56505 50331 56563 50337
rect 57054 50328 57060 50340
rect 57112 50328 57118 50380
rect 57882 50368 57888 50380
rect 57843 50340 57888 50368
rect 57882 50328 57888 50340
rect 57940 50328 57946 50380
rect 29822 50300 29828 50312
rect 29783 50272 29828 50300
rect 29822 50260 29828 50272
rect 29880 50260 29886 50312
rect 29917 50303 29975 50309
rect 29917 50269 29929 50303
rect 29963 50269 29975 50303
rect 29917 50263 29975 50269
rect 27930 50204 28948 50232
rect 27930 50201 27942 50204
rect 27884 50195 27942 50201
rect 29932 50176 29960 50263
rect 30006 50260 30012 50312
rect 30064 50300 30070 50312
rect 30193 50303 30251 50309
rect 30064 50272 30157 50300
rect 30064 50260 30070 50272
rect 30193 50269 30205 50303
rect 30239 50300 30251 50303
rect 30282 50300 30288 50312
rect 30239 50272 30288 50300
rect 30239 50269 30251 50272
rect 30193 50263 30251 50269
rect 30282 50260 30288 50272
rect 30340 50260 30346 50312
rect 30926 50300 30932 50312
rect 30887 50272 30932 50300
rect 30926 50260 30932 50272
rect 30984 50260 30990 50312
rect 31021 50303 31079 50309
rect 31021 50269 31033 50303
rect 31067 50269 31079 50303
rect 32122 50300 32128 50312
rect 32083 50272 32128 50300
rect 31021 50263 31079 50269
rect 30098 50192 30104 50244
rect 30156 50232 30162 50244
rect 31036 50232 31064 50263
rect 32122 50260 32128 50272
rect 32180 50260 32186 50312
rect 30156 50204 31064 50232
rect 32392 50235 32450 50241
rect 30156 50192 30162 50204
rect 32392 50201 32404 50235
rect 32438 50232 32450 50235
rect 33134 50232 33140 50244
rect 32438 50204 33140 50232
rect 32438 50201 32450 50204
rect 32392 50195 32450 50201
rect 33134 50192 33140 50204
rect 33192 50192 33198 50244
rect 18509 50167 18567 50173
rect 18509 50133 18521 50167
rect 18555 50133 18567 50167
rect 20622 50164 20628 50176
rect 20583 50136 20628 50164
rect 18509 50127 18567 50133
rect 20622 50124 20628 50136
rect 20680 50124 20686 50176
rect 22186 50164 22192 50176
rect 22147 50136 22192 50164
rect 22186 50124 22192 50136
rect 22244 50124 22250 50176
rect 29914 50124 29920 50176
rect 29972 50124 29978 50176
rect 32306 50124 32312 50176
rect 32364 50164 32370 50176
rect 33962 50164 33968 50176
rect 32364 50136 33968 50164
rect 32364 50124 32370 50136
rect 33962 50124 33968 50136
rect 34020 50124 34026 50176
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 18785 49963 18843 49969
rect 18785 49929 18797 49963
rect 18831 49960 18843 49963
rect 19426 49960 19432 49972
rect 18831 49932 19432 49960
rect 18831 49929 18843 49932
rect 18785 49923 18843 49929
rect 19426 49920 19432 49932
rect 19484 49920 19490 49972
rect 19978 49920 19984 49972
rect 20036 49960 20042 49972
rect 20441 49963 20499 49969
rect 20441 49960 20453 49963
rect 20036 49932 20453 49960
rect 20036 49920 20042 49932
rect 20441 49929 20453 49932
rect 20487 49929 20499 49963
rect 20622 49960 20628 49972
rect 20583 49932 20628 49960
rect 20441 49923 20499 49929
rect 20622 49920 20628 49932
rect 20680 49920 20686 49972
rect 29546 49920 29552 49972
rect 29604 49960 29610 49972
rect 29641 49963 29699 49969
rect 29641 49960 29653 49963
rect 29604 49932 29653 49960
rect 29604 49920 29610 49932
rect 29641 49929 29653 49932
rect 29687 49960 29699 49963
rect 30098 49960 30104 49972
rect 29687 49932 30104 49960
rect 29687 49929 29699 49932
rect 29641 49923 29699 49929
rect 30098 49920 30104 49932
rect 30156 49920 30162 49972
rect 30926 49960 30932 49972
rect 30839 49932 30932 49960
rect 30926 49920 30932 49932
rect 30984 49920 30990 49972
rect 32306 49960 32312 49972
rect 32267 49932 32312 49960
rect 32306 49920 32312 49932
rect 32364 49920 32370 49972
rect 32490 49960 32496 49972
rect 32451 49932 32496 49960
rect 32490 49920 32496 49932
rect 32548 49920 32554 49972
rect 32674 49960 32680 49972
rect 32635 49932 32680 49960
rect 32674 49920 32680 49932
rect 32732 49920 32738 49972
rect 33134 49960 33140 49972
rect 33095 49932 33140 49960
rect 33134 49920 33140 49932
rect 33192 49920 33198 49972
rect 19797 49895 19855 49901
rect 19797 49892 19809 49895
rect 18984 49864 19809 49892
rect 18984 49833 19012 49864
rect 19797 49861 19809 49864
rect 19843 49861 19855 49895
rect 20254 49892 20260 49904
rect 20215 49864 20260 49892
rect 19797 49855 19855 49861
rect 20254 49852 20260 49864
rect 20312 49852 20318 49904
rect 24026 49852 24032 49904
rect 24084 49892 24090 49904
rect 24489 49895 24547 49901
rect 24489 49892 24501 49895
rect 24084 49864 24501 49892
rect 24084 49852 24090 49864
rect 24489 49861 24501 49864
rect 24535 49861 24547 49895
rect 27614 49892 27620 49904
rect 27575 49864 27620 49892
rect 24489 49855 24547 49861
rect 27614 49852 27620 49864
rect 27672 49892 27678 49904
rect 28528 49895 28586 49901
rect 27672 49864 28488 49892
rect 27672 49852 27678 49864
rect 18969 49827 19027 49833
rect 18969 49793 18981 49827
rect 19015 49793 19027 49827
rect 18969 49787 19027 49793
rect 19613 49827 19671 49833
rect 19613 49793 19625 49827
rect 19659 49824 19671 49827
rect 20070 49824 20076 49836
rect 19659 49796 20076 49824
rect 19659 49793 19671 49796
rect 19613 49787 19671 49793
rect 20070 49784 20076 49796
rect 20128 49784 20134 49836
rect 20530 49824 20536 49836
rect 20491 49796 20536 49824
rect 20530 49784 20536 49796
rect 20588 49784 20594 49836
rect 22649 49827 22707 49833
rect 22649 49793 22661 49827
rect 22695 49824 22707 49827
rect 22695 49796 23428 49824
rect 22695 49793 22707 49796
rect 22649 49787 22707 49793
rect 3418 49716 3424 49768
rect 3476 49756 3482 49768
rect 9674 49756 9680 49768
rect 3476 49728 9680 49756
rect 3476 49716 3482 49728
rect 9674 49716 9680 49728
rect 9732 49716 9738 49768
rect 19429 49759 19487 49765
rect 19429 49725 19441 49759
rect 19475 49756 19487 49759
rect 20162 49756 20168 49768
rect 19475 49728 20168 49756
rect 19475 49725 19487 49728
rect 19429 49719 19487 49725
rect 20162 49716 20168 49728
rect 20220 49756 20226 49768
rect 20622 49756 20628 49768
rect 20220 49728 20628 49756
rect 20220 49716 20226 49728
rect 20622 49716 20628 49728
rect 20680 49716 20686 49768
rect 20809 49759 20867 49765
rect 20809 49725 20821 49759
rect 20855 49756 20867 49759
rect 22002 49756 22008 49768
rect 20855 49728 22008 49756
rect 20855 49725 20867 49728
rect 20809 49719 20867 49725
rect 22002 49716 22008 49728
rect 22060 49716 22066 49768
rect 23293 49759 23351 49765
rect 23293 49725 23305 49759
rect 23339 49725 23351 49759
rect 23400 49756 23428 49796
rect 23474 49784 23480 49836
rect 23532 49824 23538 49836
rect 23532 49796 23577 49824
rect 23532 49784 23538 49796
rect 24118 49784 24124 49836
rect 24176 49824 24182 49836
rect 24305 49827 24363 49833
rect 24305 49824 24317 49827
rect 24176 49796 24317 49824
rect 24176 49784 24182 49796
rect 24305 49793 24317 49796
rect 24351 49793 24363 49827
rect 24305 49787 24363 49793
rect 24394 49784 24400 49836
rect 24452 49824 24458 49836
rect 27433 49827 27491 49833
rect 27433 49824 27445 49827
rect 24452 49796 24497 49824
rect 25608 49796 27445 49824
rect 24452 49784 24458 49796
rect 25608 49768 25636 49796
rect 27433 49793 27445 49796
rect 27479 49793 27491 49827
rect 28258 49824 28264 49836
rect 28219 49796 28264 49824
rect 27433 49787 27491 49793
rect 28258 49784 28264 49796
rect 28316 49784 28322 49836
rect 28460 49824 28488 49864
rect 28528 49861 28540 49895
rect 28574 49892 28586 49895
rect 30944 49892 30972 49920
rect 28574 49864 30972 49892
rect 28574 49861 28586 49864
rect 28528 49855 28586 49861
rect 31662 49852 31668 49904
rect 31720 49892 31726 49904
rect 32125 49895 32183 49901
rect 32125 49892 32137 49895
rect 31720 49864 32137 49892
rect 31720 49852 31726 49864
rect 32125 49861 32137 49864
rect 32171 49861 32183 49895
rect 32125 49855 32183 49861
rect 32401 49895 32459 49901
rect 32401 49861 32413 49895
rect 32447 49892 32459 49895
rect 33502 49892 33508 49904
rect 32447 49864 33508 49892
rect 32447 49861 32459 49864
rect 32401 49855 32459 49861
rect 33502 49852 33508 49864
rect 33560 49852 33566 49904
rect 29086 49824 29092 49836
rect 28460 49796 29092 49824
rect 29086 49784 29092 49796
rect 29144 49784 29150 49836
rect 29270 49784 29276 49836
rect 29328 49824 29334 49836
rect 30285 49827 30343 49833
rect 30285 49824 30297 49827
rect 29328 49796 30297 49824
rect 29328 49784 29334 49796
rect 30285 49793 30297 49796
rect 30331 49793 30343 49827
rect 30285 49787 30343 49793
rect 30469 49827 30527 49833
rect 30469 49793 30481 49827
rect 30515 49824 30527 49827
rect 31113 49827 31171 49833
rect 31113 49824 31125 49827
rect 30515 49796 31125 49824
rect 30515 49793 30527 49796
rect 30469 49787 30527 49793
rect 31113 49793 31125 49796
rect 31159 49793 31171 49827
rect 31113 49787 31171 49793
rect 33042 49784 33048 49836
rect 33100 49824 33106 49836
rect 37826 49833 37832 49836
rect 33321 49827 33379 49833
rect 33321 49824 33333 49827
rect 33100 49796 33333 49824
rect 33100 49784 33106 49796
rect 33321 49793 33333 49796
rect 33367 49793 33379 49827
rect 33321 49787 33379 49793
rect 37820 49787 37832 49833
rect 37884 49824 37890 49836
rect 37884 49796 37920 49824
rect 37826 49784 37832 49787
rect 37884 49784 37890 49796
rect 39206 49784 39212 49836
rect 39264 49824 39270 49836
rect 39485 49827 39543 49833
rect 39485 49824 39497 49827
rect 39264 49796 39497 49824
rect 39264 49784 39270 49796
rect 39485 49793 39497 49796
rect 39531 49824 39543 49827
rect 39942 49824 39948 49836
rect 39531 49796 39948 49824
rect 39531 49793 39543 49796
rect 39485 49787 39543 49793
rect 39942 49784 39948 49796
rect 40000 49824 40006 49836
rect 40129 49827 40187 49833
rect 40129 49824 40141 49827
rect 40000 49796 40141 49824
rect 40000 49784 40006 49796
rect 40129 49793 40141 49796
rect 40175 49793 40187 49827
rect 40310 49824 40316 49836
rect 40271 49796 40316 49824
rect 40129 49787 40187 49793
rect 40310 49784 40316 49796
rect 40368 49784 40374 49836
rect 23566 49756 23572 49768
rect 23400 49728 23572 49756
rect 23293 49719 23351 49725
rect 23308 49688 23336 49719
rect 23566 49716 23572 49728
rect 23624 49716 23630 49768
rect 23661 49759 23719 49765
rect 23661 49725 23673 49759
rect 23707 49756 23719 49759
rect 23842 49756 23848 49768
rect 23707 49728 23848 49756
rect 23707 49725 23719 49728
rect 23661 49719 23719 49725
rect 23842 49716 23848 49728
rect 23900 49716 23906 49768
rect 24670 49756 24676 49768
rect 24631 49728 24676 49756
rect 24670 49716 24676 49728
rect 24728 49716 24734 49768
rect 25409 49759 25467 49765
rect 25409 49725 25421 49759
rect 25455 49756 25467 49759
rect 25590 49756 25596 49768
rect 25455 49728 25596 49756
rect 25455 49725 25467 49728
rect 25409 49719 25467 49725
rect 25590 49716 25596 49728
rect 25648 49716 25654 49768
rect 25685 49759 25743 49765
rect 25685 49725 25697 49759
rect 25731 49756 25743 49759
rect 25774 49756 25780 49768
rect 25731 49728 25780 49756
rect 25731 49725 25743 49728
rect 25685 49719 25743 49725
rect 25774 49716 25780 49728
rect 25832 49716 25838 49768
rect 30098 49756 30104 49768
rect 30059 49728 30104 49756
rect 30098 49716 30104 49728
rect 30156 49716 30162 49768
rect 37366 49716 37372 49768
rect 37424 49756 37430 49768
rect 37553 49759 37611 49765
rect 37553 49756 37565 49759
rect 37424 49728 37565 49756
rect 37424 49716 37430 49728
rect 37553 49725 37565 49728
rect 37599 49725 37611 49759
rect 39666 49756 39672 49768
rect 39627 49728 39672 49756
rect 37553 49719 37611 49725
rect 39666 49716 39672 49728
rect 39724 49716 39730 49768
rect 40497 49759 40555 49765
rect 40497 49725 40509 49759
rect 40543 49756 40555 49759
rect 41506 49756 41512 49768
rect 40543 49728 41512 49756
rect 40543 49725 40555 49728
rect 40497 49719 40555 49725
rect 41506 49716 41512 49728
rect 41564 49716 41570 49768
rect 23474 49688 23480 49700
rect 23308 49660 23480 49688
rect 23474 49648 23480 49660
rect 23532 49688 23538 49700
rect 24121 49691 24179 49697
rect 24121 49688 24133 49691
rect 23532 49660 24133 49688
rect 23532 49648 23538 49660
rect 24121 49657 24133 49660
rect 24167 49657 24179 49691
rect 24121 49651 24179 49657
rect 22370 49580 22376 49632
rect 22428 49620 22434 49632
rect 22465 49623 22523 49629
rect 22465 49620 22477 49623
rect 22428 49592 22477 49620
rect 22428 49580 22434 49592
rect 22465 49589 22477 49592
rect 22511 49589 22523 49623
rect 38930 49620 38936 49632
rect 38891 49592 38936 49620
rect 22465 49583 22523 49589
rect 38930 49580 38936 49592
rect 38988 49580 38994 49632
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 19242 49376 19248 49428
rect 19300 49416 19306 49428
rect 19300 49388 20300 49416
rect 19300 49376 19306 49388
rect 19242 49280 19248 49292
rect 19203 49252 19248 49280
rect 19242 49240 19248 49252
rect 19300 49240 19306 49292
rect 19512 49215 19570 49221
rect 19512 49181 19524 49215
rect 19558 49181 19570 49215
rect 20272 49212 20300 49388
rect 23566 49376 23572 49428
rect 23624 49416 23630 49428
rect 23845 49419 23903 49425
rect 23845 49416 23857 49419
rect 23624 49388 23857 49416
rect 23624 49376 23630 49388
rect 23845 49385 23857 49388
rect 23891 49385 23903 49419
rect 23845 49379 23903 49385
rect 29178 49376 29184 49428
rect 29236 49416 29242 49428
rect 29454 49416 29460 49428
rect 29236 49388 29460 49416
rect 29236 49376 29242 49388
rect 29454 49376 29460 49388
rect 29512 49416 29518 49428
rect 29549 49419 29607 49425
rect 29549 49416 29561 49419
rect 29512 49388 29561 49416
rect 29512 49376 29518 49388
rect 29549 49385 29561 49388
rect 29595 49385 29607 49419
rect 29549 49379 29607 49385
rect 29914 49376 29920 49428
rect 29972 49416 29978 49428
rect 30009 49419 30067 49425
rect 30009 49416 30021 49419
rect 29972 49388 30021 49416
rect 29972 49376 29978 49388
rect 30009 49385 30021 49388
rect 30055 49385 30067 49419
rect 30009 49379 30067 49385
rect 39942 49376 39948 49428
rect 40000 49416 40006 49428
rect 41233 49419 41291 49425
rect 41233 49416 41245 49419
rect 40000 49388 41245 49416
rect 40000 49376 40006 49388
rect 41233 49385 41245 49388
rect 41279 49385 41291 49419
rect 41233 49379 41291 49385
rect 23017 49351 23075 49357
rect 23017 49317 23029 49351
rect 23063 49348 23075 49351
rect 28997 49351 29055 49357
rect 23063 49320 23520 49348
rect 23063 49317 23075 49320
rect 23017 49311 23075 49317
rect 23492 49289 23520 49320
rect 28997 49317 29009 49351
rect 29043 49348 29055 49351
rect 29043 49320 29868 49348
rect 29043 49317 29055 49320
rect 28997 49311 29055 49317
rect 23477 49283 23535 49289
rect 23477 49249 23489 49283
rect 23523 49280 23535 49283
rect 24118 49280 24124 49292
rect 23523 49252 24124 49280
rect 23523 49249 23535 49252
rect 23477 49243 23535 49249
rect 24118 49240 24124 49252
rect 24176 49240 24182 49292
rect 26050 49240 26056 49292
rect 26108 49280 26114 49292
rect 29730 49280 29736 49292
rect 26108 49252 26464 49280
rect 29691 49252 29736 49280
rect 26108 49240 26114 49252
rect 21634 49212 21640 49224
rect 20272 49184 21640 49212
rect 19512 49175 19570 49181
rect 19426 49104 19432 49156
rect 19484 49144 19490 49156
rect 19536 49144 19564 49175
rect 21634 49172 21640 49184
rect 21692 49172 21698 49224
rect 21904 49215 21962 49221
rect 21904 49181 21916 49215
rect 21950 49212 21962 49215
rect 22186 49212 22192 49224
rect 21950 49184 22192 49212
rect 21950 49181 21962 49184
rect 21904 49175 21962 49181
rect 22186 49172 22192 49184
rect 22244 49172 22250 49224
rect 23658 49212 23664 49224
rect 23619 49184 23664 49212
rect 23658 49172 23664 49184
rect 23716 49172 23722 49224
rect 24397 49215 24455 49221
rect 24397 49181 24409 49215
rect 24443 49212 24455 49215
rect 25038 49212 25044 49224
rect 24443 49184 25044 49212
rect 24443 49181 24455 49184
rect 24397 49175 24455 49181
rect 25038 49172 25044 49184
rect 25096 49172 25102 49224
rect 26436 49221 26464 49252
rect 29730 49240 29736 49252
rect 29788 49240 29794 49292
rect 26237 49215 26295 49221
rect 26237 49212 26249 49215
rect 25792 49184 26249 49212
rect 19484 49116 19564 49144
rect 19484 49104 19490 49116
rect 23750 49104 23756 49156
rect 23808 49144 23814 49156
rect 24642 49147 24700 49153
rect 24642 49144 24654 49147
rect 23808 49116 24654 49144
rect 23808 49104 23814 49116
rect 24642 49113 24654 49116
rect 24688 49113 24700 49147
rect 24642 49107 24700 49113
rect 20622 49076 20628 49088
rect 20583 49048 20628 49076
rect 20622 49036 20628 49048
rect 20680 49036 20686 49088
rect 24026 49036 24032 49088
rect 24084 49076 24090 49088
rect 25792 49085 25820 49184
rect 26237 49181 26249 49184
rect 26283 49181 26295 49215
rect 26237 49175 26295 49181
rect 26421 49215 26479 49221
rect 26421 49181 26433 49215
rect 26467 49181 26479 49215
rect 26421 49175 26479 49181
rect 27617 49215 27675 49221
rect 27617 49181 27629 49215
rect 27663 49212 27675 49215
rect 28258 49212 28264 49224
rect 27663 49184 28264 49212
rect 27663 49181 27675 49184
rect 27617 49175 27675 49181
rect 28258 49172 28264 49184
rect 28316 49172 28322 49224
rect 29546 49212 29552 49224
rect 29507 49184 29552 49212
rect 29546 49172 29552 49184
rect 29604 49172 29610 49224
rect 29840 49221 29868 49320
rect 38930 49240 38936 49292
rect 38988 49280 38994 49292
rect 39850 49280 39856 49292
rect 38988 49252 39856 49280
rect 38988 49240 38994 49252
rect 39850 49240 39856 49252
rect 39908 49240 39914 49292
rect 48958 49280 48964 49292
rect 42076 49252 43116 49280
rect 48919 49252 48964 49280
rect 29825 49215 29883 49221
rect 29825 49181 29837 49215
rect 29871 49212 29883 49215
rect 30098 49212 30104 49224
rect 29871 49184 30104 49212
rect 29871 49181 29883 49184
rect 29825 49175 29883 49181
rect 30098 49172 30104 49184
rect 30156 49172 30162 49224
rect 30745 49215 30803 49221
rect 30745 49181 30757 49215
rect 30791 49212 30803 49215
rect 32122 49212 32128 49224
rect 30791 49184 32128 49212
rect 30791 49181 30803 49184
rect 30745 49175 30803 49181
rect 32122 49172 32128 49184
rect 32180 49212 32186 49224
rect 34701 49215 34759 49221
rect 34701 49212 34713 49215
rect 32180 49184 34713 49212
rect 32180 49172 32186 49184
rect 34701 49181 34713 49184
rect 34747 49212 34759 49215
rect 37366 49212 37372 49224
rect 34747 49184 37372 49212
rect 34747 49181 34759 49184
rect 34701 49175 34759 49181
rect 37366 49172 37372 49184
rect 37424 49172 37430 49224
rect 40126 49212 40132 49224
rect 40087 49184 40132 49212
rect 40126 49172 40132 49184
rect 40184 49212 40190 49224
rect 40310 49212 40316 49224
rect 40184 49184 40316 49212
rect 40184 49172 40190 49184
rect 40310 49172 40316 49184
rect 40368 49212 40374 49224
rect 41141 49215 41199 49221
rect 41141 49212 41153 49215
rect 40368 49184 41153 49212
rect 40368 49172 40374 49184
rect 41141 49181 41153 49184
rect 41187 49181 41199 49215
rect 41141 49175 41199 49181
rect 41782 49172 41788 49224
rect 41840 49212 41846 49224
rect 42076 49221 42104 49252
rect 42061 49215 42119 49221
rect 42061 49212 42073 49215
rect 41840 49184 42073 49212
rect 41840 49172 41846 49184
rect 42061 49181 42073 49184
rect 42107 49181 42119 49215
rect 42702 49212 42708 49224
rect 42061 49175 42119 49181
rect 42260 49184 42708 49212
rect 27890 49153 27896 49156
rect 27884 49107 27896 49153
rect 27948 49144 27954 49156
rect 30558 49144 30564 49156
rect 27948 49116 27984 49144
rect 30519 49116 30564 49144
rect 27890 49104 27896 49107
rect 27948 49104 27954 49116
rect 30558 49104 30564 49116
rect 30616 49104 30622 49156
rect 34238 49104 34244 49156
rect 34296 49144 34302 49156
rect 34946 49147 35004 49153
rect 34946 49144 34958 49147
rect 34296 49116 34958 49144
rect 34296 49104 34302 49116
rect 34946 49113 34958 49116
rect 34992 49113 35004 49147
rect 34946 49107 35004 49113
rect 37274 49104 37280 49156
rect 37332 49144 37338 49156
rect 37614 49147 37672 49153
rect 37614 49144 37626 49147
rect 37332 49116 37626 49144
rect 37332 49104 37338 49116
rect 37614 49113 37626 49116
rect 37660 49113 37672 49147
rect 37614 49107 37672 49113
rect 41966 49104 41972 49156
rect 42024 49144 42030 49156
rect 42260 49153 42288 49184
rect 42702 49172 42708 49184
rect 42760 49212 42766 49224
rect 43088 49221 43116 49252
rect 48958 49240 48964 49252
rect 49016 49240 49022 49292
rect 42889 49215 42947 49221
rect 42889 49212 42901 49215
rect 42760 49184 42901 49212
rect 42760 49172 42766 49184
rect 42889 49181 42901 49184
rect 42935 49181 42947 49215
rect 42889 49175 42947 49181
rect 43073 49215 43131 49221
rect 43073 49181 43085 49215
rect 43119 49181 43131 49215
rect 47762 49212 47768 49224
rect 47723 49184 47768 49212
rect 43073 49175 43131 49181
rect 47762 49172 47768 49184
rect 47820 49172 47826 49224
rect 56594 49172 56600 49224
rect 56652 49212 56658 49224
rect 57057 49215 57115 49221
rect 57057 49212 57069 49215
rect 56652 49184 57069 49212
rect 56652 49172 56658 49184
rect 57057 49181 57069 49184
rect 57103 49181 57115 49215
rect 57057 49175 57115 49181
rect 42245 49147 42303 49153
rect 42245 49144 42257 49147
rect 42024 49116 42257 49144
rect 42024 49104 42030 49116
rect 42245 49113 42257 49116
rect 42291 49113 42303 49147
rect 42245 49107 42303 49113
rect 42429 49147 42487 49153
rect 42429 49113 42441 49147
rect 42475 49144 42487 49147
rect 43530 49144 43536 49156
rect 42475 49116 43536 49144
rect 42475 49113 42487 49116
rect 42429 49107 42487 49113
rect 43530 49104 43536 49116
rect 43588 49104 43594 49156
rect 47949 49147 48007 49153
rect 47949 49113 47961 49147
rect 47995 49144 48007 49147
rect 48222 49144 48228 49156
rect 47995 49116 48228 49144
rect 47995 49113 48007 49116
rect 47949 49107 48007 49113
rect 48222 49104 48228 49116
rect 48280 49104 48286 49156
rect 57072 49144 57100 49175
rect 57238 49172 57244 49224
rect 57296 49212 57302 49224
rect 57885 49215 57943 49221
rect 57885 49212 57897 49215
rect 57296 49184 57897 49212
rect 57296 49172 57302 49184
rect 57885 49181 57897 49184
rect 57931 49181 57943 49215
rect 57885 49175 57943 49181
rect 57606 49144 57612 49156
rect 57072 49116 57612 49144
rect 57606 49104 57612 49116
rect 57664 49104 57670 49156
rect 25777 49079 25835 49085
rect 25777 49076 25789 49079
rect 24084 49048 25789 49076
rect 24084 49036 24090 49048
rect 25777 49045 25789 49048
rect 25823 49045 25835 49079
rect 25777 49039 25835 49045
rect 26605 49079 26663 49085
rect 26605 49045 26617 49079
rect 26651 49076 26663 49079
rect 27154 49076 27160 49088
rect 26651 49048 27160 49076
rect 26651 49045 26663 49048
rect 26605 49039 26663 49045
rect 27154 49036 27160 49048
rect 27212 49036 27218 49088
rect 36078 49076 36084 49088
rect 36039 49048 36084 49076
rect 36078 49036 36084 49048
rect 36136 49036 36142 49088
rect 38746 49076 38752 49088
rect 38707 49048 38752 49076
rect 38746 49036 38752 49048
rect 38804 49036 38810 49088
rect 41601 49079 41659 49085
rect 41601 49045 41613 49079
rect 41647 49076 41659 49079
rect 42886 49076 42892 49088
rect 41647 49048 42892 49076
rect 41647 49045 41659 49048
rect 41601 49039 41659 49045
rect 42886 49036 42892 49048
rect 42944 49036 42950 49088
rect 43165 49079 43223 49085
rect 43165 49045 43177 49079
rect 43211 49076 43223 49079
rect 44450 49076 44456 49088
rect 43211 49048 44456 49076
rect 43211 49045 43223 49048
rect 43165 49039 43223 49045
rect 44450 49036 44456 49048
rect 44508 49036 44514 49088
rect 57146 49076 57152 49088
rect 57107 49048 57152 49076
rect 57146 49036 57152 49048
rect 57204 49036 57210 49088
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 23474 48872 23480 48884
rect 23435 48844 23480 48872
rect 23474 48832 23480 48844
rect 23532 48872 23538 48884
rect 24302 48872 24308 48884
rect 23532 48844 24308 48872
rect 23532 48832 23538 48844
rect 24302 48832 24308 48844
rect 24360 48832 24366 48884
rect 26973 48875 27031 48881
rect 26973 48841 26985 48875
rect 27019 48841 27031 48875
rect 26973 48835 27031 48841
rect 27801 48875 27859 48881
rect 27801 48841 27813 48875
rect 27847 48872 27859 48875
rect 27890 48872 27896 48884
rect 27847 48844 27896 48872
rect 27847 48841 27859 48844
rect 27801 48835 27859 48841
rect 19150 48804 19156 48816
rect 7852 48776 19156 48804
rect 7852 48745 7880 48776
rect 19150 48764 19156 48776
rect 19208 48764 19214 48816
rect 20162 48804 20168 48816
rect 20123 48776 20168 48804
rect 20162 48764 20168 48776
rect 20220 48764 20226 48816
rect 20254 48764 20260 48816
rect 20312 48804 20318 48816
rect 20312 48776 20484 48804
rect 20312 48764 20318 48776
rect 20456 48745 20484 48776
rect 21634 48764 21640 48816
rect 21692 48804 21698 48816
rect 25308 48807 25366 48813
rect 21692 48776 25084 48804
rect 21692 48764 21698 48776
rect 22112 48745 22140 48776
rect 25056 48748 25084 48776
rect 25308 48773 25320 48807
rect 25354 48804 25366 48807
rect 26988 48804 27016 48835
rect 27890 48832 27896 48844
rect 27948 48832 27954 48884
rect 34238 48872 34244 48884
rect 34199 48844 34244 48872
rect 34238 48832 34244 48844
rect 34296 48832 34302 48884
rect 36078 48832 36084 48884
rect 36136 48872 36142 48884
rect 47762 48872 47768 48884
rect 36136 48844 47768 48872
rect 36136 48832 36142 48844
rect 47762 48832 47768 48844
rect 47820 48832 47826 48884
rect 48222 48872 48228 48884
rect 48183 48844 48228 48872
rect 48222 48832 48228 48844
rect 48280 48832 48286 48884
rect 28813 48807 28871 48813
rect 28813 48804 28825 48807
rect 25354 48776 27016 48804
rect 28000 48776 28825 48804
rect 25354 48773 25366 48776
rect 25308 48767 25366 48773
rect 22370 48745 22376 48748
rect 7837 48739 7895 48745
rect 7837 48705 7849 48739
rect 7883 48705 7895 48739
rect 7837 48699 7895 48705
rect 20441 48739 20499 48745
rect 20441 48705 20453 48739
rect 20487 48705 20499 48739
rect 20441 48699 20499 48705
rect 22097 48739 22155 48745
rect 22097 48705 22109 48739
rect 22143 48736 22155 48739
rect 22364 48736 22376 48745
rect 22143 48708 22177 48736
rect 22331 48708 22376 48736
rect 22143 48705 22155 48708
rect 22097 48699 22155 48705
rect 22364 48699 22376 48708
rect 22370 48696 22376 48699
rect 22428 48696 22434 48748
rect 24026 48736 24032 48748
rect 23987 48708 24032 48736
rect 24026 48696 24032 48708
rect 24084 48696 24090 48748
rect 24302 48736 24308 48748
rect 24263 48708 24308 48736
rect 24302 48696 24308 48708
rect 24360 48696 24366 48748
rect 25038 48736 25044 48748
rect 24999 48708 25044 48736
rect 25038 48696 25044 48708
rect 25096 48696 25102 48748
rect 27154 48736 27160 48748
rect 27115 48708 27160 48736
rect 27154 48696 27160 48708
rect 27212 48696 27218 48748
rect 28000 48745 28028 48776
rect 28813 48773 28825 48776
rect 28859 48773 28871 48807
rect 29362 48804 29368 48816
rect 28813 48767 28871 48773
rect 28966 48776 29368 48804
rect 27985 48739 28043 48745
rect 27985 48705 27997 48739
rect 28031 48705 28043 48739
rect 27985 48699 28043 48705
rect 28074 48696 28080 48748
rect 28132 48736 28138 48748
rect 28629 48739 28687 48745
rect 28629 48736 28641 48739
rect 28132 48708 28641 48736
rect 28132 48696 28138 48708
rect 28629 48705 28641 48708
rect 28675 48736 28687 48739
rect 28966 48736 28994 48776
rect 29362 48764 29368 48776
rect 29420 48764 29426 48816
rect 29638 48764 29644 48816
rect 29696 48804 29702 48816
rect 29696 48776 29741 48804
rect 29696 48764 29702 48776
rect 31938 48764 31944 48816
rect 31996 48804 32002 48816
rect 33873 48807 33931 48813
rect 33873 48804 33885 48807
rect 31996 48776 33885 48804
rect 31996 48764 32002 48776
rect 33873 48773 33885 48776
rect 33919 48773 33931 48807
rect 33873 48767 33931 48773
rect 33965 48807 34023 48813
rect 33965 48773 33977 48807
rect 34011 48804 34023 48807
rect 36096 48804 36124 48832
rect 41782 48804 41788 48816
rect 34011 48776 36124 48804
rect 41743 48776 41788 48804
rect 34011 48773 34023 48776
rect 33965 48767 34023 48773
rect 41782 48764 41788 48776
rect 41840 48764 41846 48816
rect 28675 48708 28994 48736
rect 28675 48705 28687 48708
rect 28629 48699 28687 48705
rect 29454 48702 29460 48754
rect 29512 48742 29518 48754
rect 29512 48714 29557 48742
rect 33686 48736 33692 48748
rect 29512 48702 29518 48714
rect 33647 48708 33692 48736
rect 33686 48696 33692 48708
rect 33744 48696 33750 48748
rect 34057 48739 34115 48745
rect 34057 48705 34069 48739
rect 34103 48705 34115 48739
rect 37366 48736 37372 48748
rect 37327 48708 37372 48736
rect 34057 48699 34115 48705
rect 8478 48668 8484 48680
rect 8439 48640 8484 48668
rect 8478 48628 8484 48640
rect 8536 48628 8542 48680
rect 8665 48671 8723 48677
rect 8665 48637 8677 48671
rect 8711 48637 8723 48671
rect 9674 48668 9680 48680
rect 9635 48640 9680 48668
rect 8665 48631 8723 48637
rect 7929 48603 7987 48609
rect 7929 48569 7941 48603
rect 7975 48600 7987 48603
rect 8680 48600 8708 48631
rect 9674 48628 9680 48640
rect 9732 48628 9738 48680
rect 19702 48628 19708 48680
rect 19760 48668 19766 48680
rect 20257 48671 20315 48677
rect 20257 48668 20269 48671
rect 19760 48640 20269 48668
rect 19760 48628 19766 48640
rect 20257 48637 20269 48640
rect 20303 48668 20315 48671
rect 20622 48668 20628 48680
rect 20303 48640 20628 48668
rect 20303 48637 20315 48640
rect 20257 48631 20315 48637
rect 20622 48628 20628 48640
rect 20680 48628 20686 48680
rect 24213 48671 24271 48677
rect 24213 48637 24225 48671
rect 24259 48668 24271 48671
rect 24394 48668 24400 48680
rect 24259 48640 24400 48668
rect 24259 48637 24271 48640
rect 24213 48631 24271 48637
rect 24394 48628 24400 48640
rect 24452 48668 24458 48680
rect 28445 48671 28503 48677
rect 24452 48640 24992 48668
rect 24452 48628 24458 48640
rect 7975 48572 8708 48600
rect 7975 48569 7987 48572
rect 7929 48563 7987 48569
rect 19978 48492 19984 48544
rect 20036 48532 20042 48544
rect 20165 48535 20223 48541
rect 20165 48532 20177 48535
rect 20036 48504 20177 48532
rect 20036 48492 20042 48504
rect 20165 48501 20177 48504
rect 20211 48501 20223 48535
rect 20165 48495 20223 48501
rect 20625 48535 20683 48541
rect 20625 48501 20637 48535
rect 20671 48532 20683 48535
rect 21358 48532 21364 48544
rect 20671 48504 21364 48532
rect 20671 48501 20683 48504
rect 20625 48495 20683 48501
rect 21358 48492 21364 48504
rect 21416 48492 21422 48544
rect 24118 48532 24124 48544
rect 24079 48504 24124 48532
rect 24118 48492 24124 48504
rect 24176 48492 24182 48544
rect 24394 48492 24400 48544
rect 24452 48532 24458 48544
rect 24489 48535 24547 48541
rect 24489 48532 24501 48535
rect 24452 48504 24501 48532
rect 24452 48492 24458 48504
rect 24489 48501 24501 48504
rect 24535 48501 24547 48535
rect 24964 48532 24992 48640
rect 28445 48637 28457 48671
rect 28491 48668 28503 48671
rect 29273 48671 29331 48677
rect 28491 48640 28994 48668
rect 28491 48637 28503 48640
rect 28445 48631 28503 48637
rect 28966 48612 28994 48640
rect 29273 48637 29285 48671
rect 29319 48637 29331 48671
rect 29273 48631 29331 48637
rect 28966 48572 29000 48612
rect 28994 48560 29000 48572
rect 29052 48600 29058 48612
rect 29178 48600 29184 48612
rect 29052 48572 29184 48600
rect 29052 48560 29058 48572
rect 29178 48560 29184 48572
rect 29236 48560 29242 48612
rect 29288 48600 29316 48631
rect 32582 48628 32588 48680
rect 32640 48668 32646 48680
rect 34072 48668 34100 48699
rect 37366 48696 37372 48708
rect 37424 48696 37430 48748
rect 37636 48739 37694 48745
rect 37636 48705 37648 48739
rect 37682 48736 37694 48739
rect 38194 48736 38200 48748
rect 37682 48708 38200 48736
rect 37682 48705 37694 48708
rect 37636 48699 37694 48705
rect 38194 48696 38200 48708
rect 38252 48696 38258 48748
rect 38746 48696 38752 48748
rect 38804 48736 38810 48748
rect 39761 48739 39819 48745
rect 39761 48736 39773 48739
rect 38804 48708 39773 48736
rect 38804 48696 38810 48708
rect 39761 48705 39773 48708
rect 39807 48736 39819 48739
rect 39942 48736 39948 48748
rect 39807 48708 39948 48736
rect 39807 48705 39819 48708
rect 39761 48699 39819 48705
rect 39942 48696 39948 48708
rect 40000 48736 40006 48748
rect 40405 48739 40463 48745
rect 40405 48736 40417 48739
rect 40000 48708 40417 48736
rect 40000 48696 40006 48708
rect 40405 48705 40417 48708
rect 40451 48705 40463 48739
rect 40405 48699 40463 48705
rect 41693 48739 41751 48745
rect 41693 48705 41705 48739
rect 41739 48705 41751 48739
rect 41874 48736 41880 48748
rect 41835 48708 41880 48736
rect 41693 48699 41751 48705
rect 39206 48668 39212 48680
rect 32640 48640 34100 48668
rect 39167 48640 39212 48668
rect 32640 48628 32646 48640
rect 39206 48628 39212 48640
rect 39264 48628 39270 48680
rect 39577 48671 39635 48677
rect 39577 48637 39589 48671
rect 39623 48637 39635 48671
rect 39577 48631 39635 48637
rect 39669 48671 39727 48677
rect 39669 48637 39681 48671
rect 39715 48668 39727 48671
rect 40126 48668 40132 48680
rect 39715 48640 40132 48668
rect 39715 48637 39727 48640
rect 39669 48631 39727 48637
rect 29546 48600 29552 48612
rect 29288 48572 29552 48600
rect 29546 48560 29552 48572
rect 29604 48560 29610 48612
rect 38749 48603 38807 48609
rect 38749 48569 38761 48603
rect 38795 48600 38807 48603
rect 39224 48600 39252 48628
rect 38795 48572 39252 48600
rect 38795 48569 38807 48572
rect 38749 48563 38807 48569
rect 26421 48535 26479 48541
rect 26421 48532 26433 48535
rect 24964 48504 26433 48532
rect 24489 48495 24547 48501
rect 26421 48501 26433 48504
rect 26467 48501 26479 48535
rect 39592 48532 39620 48631
rect 40126 48628 40132 48640
rect 40184 48668 40190 48680
rect 40586 48668 40592 48680
rect 40184 48640 40592 48668
rect 40184 48628 40190 48640
rect 40586 48628 40592 48640
rect 40644 48628 40650 48680
rect 40681 48671 40739 48677
rect 40681 48637 40693 48671
rect 40727 48668 40739 48671
rect 41138 48668 41144 48680
rect 40727 48640 41144 48668
rect 40727 48637 40739 48640
rect 40681 48631 40739 48637
rect 41138 48628 41144 48640
rect 41196 48668 41202 48680
rect 41708 48668 41736 48699
rect 41874 48696 41880 48708
rect 41932 48696 41938 48748
rect 42429 48739 42487 48745
rect 42429 48705 42441 48739
rect 42475 48736 42487 48739
rect 43625 48739 43683 48745
rect 43625 48736 43637 48739
rect 42475 48708 43637 48736
rect 42475 48705 42487 48708
rect 42429 48699 42487 48705
rect 43625 48705 43637 48708
rect 43671 48705 43683 48739
rect 43625 48699 43683 48705
rect 43809 48739 43867 48745
rect 43809 48705 43821 48739
rect 43855 48705 43867 48739
rect 43809 48699 43867 48705
rect 44729 48739 44787 48745
rect 44729 48705 44741 48739
rect 44775 48705 44787 48739
rect 44910 48736 44916 48748
rect 44871 48708 44916 48736
rect 44729 48699 44787 48705
rect 42444 48668 42472 48699
rect 41196 48640 42472 48668
rect 41196 48628 41202 48640
rect 42518 48628 42524 48680
rect 42576 48668 42582 48680
rect 42613 48671 42671 48677
rect 42613 48668 42625 48671
rect 42576 48640 42625 48668
rect 42576 48628 42582 48640
rect 42613 48637 42625 48640
rect 42659 48637 42671 48671
rect 42613 48631 42671 48637
rect 42702 48628 42708 48680
rect 42760 48668 42766 48680
rect 42889 48671 42947 48677
rect 42889 48668 42901 48671
rect 42760 48640 42901 48668
rect 42760 48628 42766 48640
rect 42889 48637 42901 48640
rect 42935 48637 42947 48671
rect 42889 48631 42947 48637
rect 42981 48671 43039 48677
rect 42981 48637 42993 48671
rect 43027 48668 43039 48671
rect 43824 48668 43852 48699
rect 43027 48640 43852 48668
rect 44744 48668 44772 48699
rect 44910 48696 44916 48708
rect 44968 48696 44974 48748
rect 45002 48696 45008 48748
rect 45060 48736 45066 48748
rect 45186 48745 45192 48748
rect 45143 48739 45192 48745
rect 45060 48708 45105 48736
rect 45060 48696 45066 48708
rect 45143 48705 45155 48739
rect 45189 48705 45192 48739
rect 45143 48699 45192 48705
rect 45186 48696 45192 48699
rect 45244 48696 45250 48748
rect 48130 48736 48136 48748
rect 48091 48708 48136 48736
rect 48130 48696 48136 48708
rect 48188 48736 48194 48748
rect 56870 48736 56876 48748
rect 48188 48708 56876 48736
rect 48188 48696 48194 48708
rect 56870 48696 56876 48708
rect 56928 48696 56934 48748
rect 46014 48668 46020 48680
rect 44744 48640 46020 48668
rect 43027 48637 43039 48640
rect 42981 48631 43039 48637
rect 41874 48560 41880 48612
rect 41932 48600 41938 48612
rect 42996 48600 43024 48631
rect 46014 48628 46020 48640
rect 46072 48628 46078 48680
rect 41932 48572 43024 48600
rect 41932 48560 41938 48572
rect 40678 48532 40684 48544
rect 39592 48504 40684 48532
rect 26421 48495 26479 48501
rect 40678 48492 40684 48504
rect 40736 48492 40742 48544
rect 43990 48532 43996 48544
rect 43951 48504 43996 48532
rect 43990 48492 43996 48504
rect 44048 48492 44054 48544
rect 45278 48532 45284 48544
rect 45239 48504 45284 48532
rect 45278 48492 45284 48504
rect 45336 48492 45342 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 23661 48331 23719 48337
rect 23661 48297 23673 48331
rect 23707 48328 23719 48331
rect 23750 48328 23756 48340
rect 23707 48300 23756 48328
rect 23707 48297 23719 48300
rect 23661 48291 23719 48297
rect 23750 48288 23756 48300
rect 23808 48288 23814 48340
rect 37274 48328 37280 48340
rect 37235 48300 37280 48328
rect 37274 48288 37280 48300
rect 37332 48288 37338 48340
rect 38194 48288 38200 48340
rect 38252 48328 38258 48340
rect 38289 48331 38347 48337
rect 38289 48328 38301 48331
rect 38252 48300 38301 48328
rect 38252 48288 38258 48300
rect 38289 48297 38301 48300
rect 38335 48297 38347 48331
rect 41874 48328 41880 48340
rect 38289 48291 38347 48297
rect 40788 48300 41880 48328
rect 26970 48220 26976 48272
rect 27028 48260 27034 48272
rect 30190 48260 30196 48272
rect 27028 48232 30196 48260
rect 27028 48220 27034 48232
rect 30190 48220 30196 48232
rect 30248 48220 30254 48272
rect 39758 48260 39764 48272
rect 36832 48232 39764 48260
rect 25590 48192 25596 48204
rect 25551 48164 25596 48192
rect 25590 48152 25596 48164
rect 25648 48152 25654 48204
rect 28074 48192 28080 48204
rect 28035 48164 28080 48192
rect 28074 48152 28080 48164
rect 28132 48152 28138 48204
rect 19702 48124 19708 48136
rect 19663 48096 19708 48124
rect 19702 48084 19708 48096
rect 19760 48084 19766 48136
rect 19797 48127 19855 48133
rect 19797 48093 19809 48127
rect 19843 48124 19855 48127
rect 19978 48124 19984 48136
rect 19843 48096 19984 48124
rect 19843 48093 19855 48096
rect 19797 48087 19855 48093
rect 19978 48084 19984 48096
rect 20036 48084 20042 48136
rect 23842 48124 23848 48136
rect 23803 48096 23848 48124
rect 23842 48084 23848 48096
rect 23900 48084 23906 48136
rect 24394 48124 24400 48136
rect 24355 48096 24400 48124
rect 24394 48084 24400 48096
rect 24452 48084 24458 48136
rect 24578 48124 24584 48136
rect 24539 48096 24584 48124
rect 24578 48084 24584 48096
rect 24636 48084 24642 48136
rect 25317 48127 25375 48133
rect 25317 48093 25329 48127
rect 25363 48124 25375 48127
rect 26142 48124 26148 48136
rect 25363 48096 26148 48124
rect 25363 48093 25375 48096
rect 25317 48087 25375 48093
rect 26142 48084 26148 48096
rect 26200 48084 26206 48136
rect 27614 48084 27620 48136
rect 27672 48124 27678 48136
rect 27801 48127 27859 48133
rect 27801 48124 27813 48127
rect 27672 48096 27813 48124
rect 27672 48084 27678 48096
rect 27801 48093 27813 48096
rect 27847 48124 27859 48127
rect 29270 48124 29276 48136
rect 27847 48096 29276 48124
rect 27847 48093 27859 48096
rect 27801 48087 27859 48093
rect 29270 48084 29276 48096
rect 29328 48084 29334 48136
rect 31018 48084 31024 48136
rect 31076 48124 31082 48136
rect 32769 48127 32827 48133
rect 32769 48124 32781 48127
rect 31076 48096 32781 48124
rect 31076 48084 31082 48096
rect 32769 48093 32781 48096
rect 32815 48124 32827 48127
rect 34146 48124 34152 48136
rect 32815 48096 34152 48124
rect 32815 48093 32827 48096
rect 32769 48087 32827 48093
rect 34146 48084 34152 48096
rect 34204 48084 34210 48136
rect 36538 48084 36544 48136
rect 36596 48124 36602 48136
rect 36725 48127 36783 48133
rect 36725 48124 36737 48127
rect 36596 48096 36737 48124
rect 36596 48084 36602 48096
rect 36725 48093 36737 48096
rect 36771 48093 36783 48127
rect 36832 48124 36860 48232
rect 39758 48220 39764 48232
rect 39816 48260 39822 48272
rect 40129 48263 40187 48269
rect 40129 48260 40141 48263
rect 39816 48232 40141 48260
rect 39816 48220 39822 48232
rect 40129 48229 40141 48232
rect 40175 48229 40187 48263
rect 40129 48223 40187 48229
rect 37108 48164 38148 48192
rect 37108 48133 37136 48164
rect 38120 48136 38148 48164
rect 37001 48127 37059 48133
rect 37001 48124 37013 48127
rect 36832 48096 37013 48124
rect 36725 48087 36783 48093
rect 37001 48093 37013 48096
rect 37047 48093 37059 48127
rect 37001 48087 37059 48093
rect 37093 48127 37151 48133
rect 37093 48093 37105 48127
rect 37139 48093 37151 48127
rect 37093 48087 37151 48093
rect 37182 48084 37188 48136
rect 37240 48124 37246 48136
rect 37737 48127 37795 48133
rect 37737 48124 37749 48127
rect 37240 48096 37749 48124
rect 37240 48084 37246 48096
rect 37737 48093 37749 48096
rect 37783 48093 37795 48127
rect 38102 48124 38108 48136
rect 38063 48096 38108 48124
rect 37737 48087 37795 48093
rect 38102 48084 38108 48096
rect 38160 48084 38166 48136
rect 39942 48124 39948 48136
rect 39903 48096 39948 48124
rect 39942 48084 39948 48096
rect 40000 48084 40006 48136
rect 40586 48124 40592 48136
rect 40547 48096 40592 48124
rect 40586 48084 40592 48096
rect 40644 48084 40650 48136
rect 40788 48133 40816 48300
rect 41874 48288 41880 48300
rect 41932 48288 41938 48340
rect 46014 48328 46020 48340
rect 45975 48300 46020 48328
rect 46014 48288 46020 48300
rect 46072 48288 46078 48340
rect 40954 48220 40960 48272
rect 41012 48260 41018 48272
rect 45278 48260 45284 48272
rect 41012 48232 45284 48260
rect 41012 48220 41018 48232
rect 45278 48220 45284 48232
rect 45336 48220 45342 48272
rect 48130 48260 48136 48272
rect 45388 48232 48136 48260
rect 41046 48192 41052 48204
rect 41007 48164 41052 48192
rect 41046 48152 41052 48164
rect 41104 48152 41110 48204
rect 41782 48152 41788 48204
rect 41840 48192 41846 48204
rect 42521 48195 42579 48201
rect 41840 48164 42288 48192
rect 41840 48152 41846 48164
rect 40773 48127 40831 48133
rect 40773 48093 40785 48127
rect 40819 48093 40831 48127
rect 41138 48124 41144 48136
rect 41099 48096 41144 48124
rect 40773 48087 40831 48093
rect 19150 48016 19156 48068
rect 19208 48056 19214 48068
rect 30466 48056 30472 48068
rect 19208 48028 30472 48056
rect 19208 48016 19214 48028
rect 30466 48016 30472 48028
rect 30524 48016 30530 48068
rect 31938 48056 31944 48068
rect 31899 48028 31944 48056
rect 31938 48016 31944 48028
rect 31996 48016 32002 48068
rect 33042 48065 33048 48068
rect 32125 48059 32183 48065
rect 32125 48025 32137 48059
rect 32171 48025 32183 48059
rect 32125 48019 32183 48025
rect 33036 48019 33048 48065
rect 33100 48056 33106 48068
rect 36909 48059 36967 48065
rect 36909 48056 36921 48059
rect 33100 48028 33136 48056
rect 33244 48028 36921 48056
rect 19981 47991 20039 47997
rect 19981 47957 19993 47991
rect 20027 47988 20039 47991
rect 20806 47988 20812 48000
rect 20027 47960 20812 47988
rect 20027 47957 20039 47960
rect 19981 47951 20039 47957
rect 20806 47948 20812 47960
rect 20864 47948 20870 48000
rect 24762 47988 24768 48000
rect 24723 47960 24768 47988
rect 24762 47948 24768 47960
rect 24820 47948 24826 48000
rect 31754 47948 31760 48000
rect 31812 47988 31818 48000
rect 32140 47988 32168 48019
rect 33042 48016 33048 48019
rect 33100 48016 33106 48028
rect 31812 47960 32168 47988
rect 32309 47991 32367 47997
rect 31812 47948 31818 47960
rect 32309 47957 32321 47991
rect 32355 47988 32367 47991
rect 33244 47988 33272 48028
rect 36909 48025 36921 48028
rect 36955 48025 36967 48059
rect 36909 48019 36967 48025
rect 37921 48059 37979 48065
rect 37921 48025 37933 48059
rect 37967 48025 37979 48059
rect 37921 48019 37979 48025
rect 38013 48059 38071 48065
rect 38013 48025 38025 48059
rect 38059 48056 38071 48059
rect 39666 48056 39672 48068
rect 38059 48028 39672 48056
rect 38059 48025 38071 48028
rect 38013 48019 38071 48025
rect 32355 47960 33272 47988
rect 32355 47957 32367 47960
rect 32309 47951 32367 47957
rect 33318 47948 33324 48000
rect 33376 47988 33382 48000
rect 33686 47988 33692 48000
rect 33376 47960 33692 47988
rect 33376 47948 33382 47960
rect 33686 47948 33692 47960
rect 33744 47988 33750 48000
rect 34149 47991 34207 47997
rect 34149 47988 34161 47991
rect 33744 47960 34161 47988
rect 33744 47948 33750 47960
rect 34149 47957 34161 47960
rect 34195 47957 34207 47991
rect 36924 47988 36952 48019
rect 37366 47988 37372 48000
rect 36924 47960 37372 47988
rect 34149 47951 34207 47957
rect 37366 47948 37372 47960
rect 37424 47988 37430 48000
rect 37936 47988 37964 48019
rect 39666 48016 39672 48028
rect 39724 48056 39730 48068
rect 40788 48056 40816 48087
rect 41138 48084 41144 48096
rect 41196 48084 41202 48136
rect 41966 48124 41972 48136
rect 41386 48096 41972 48124
rect 39724 48028 40816 48056
rect 39724 48016 39730 48028
rect 40862 48016 40868 48068
rect 40920 48056 40926 48068
rect 41386 48056 41414 48096
rect 41966 48084 41972 48096
rect 42024 48124 42030 48136
rect 42260 48133 42288 48164
rect 42521 48161 42533 48195
rect 42567 48192 42579 48195
rect 44082 48192 44088 48204
rect 42567 48164 44088 48192
rect 42567 48161 42579 48164
rect 42521 48155 42579 48161
rect 44082 48152 44088 48164
rect 44140 48152 44146 48204
rect 44266 48152 44272 48204
rect 44324 48192 44330 48204
rect 45388 48192 45416 48232
rect 48130 48220 48136 48232
rect 48188 48220 48194 48272
rect 57238 48260 57244 48272
rect 56336 48232 57244 48260
rect 44324 48164 45416 48192
rect 45465 48195 45523 48201
rect 44324 48152 44330 48164
rect 45465 48161 45477 48195
rect 45511 48161 45523 48195
rect 45465 48155 45523 48161
rect 42061 48127 42119 48133
rect 42061 48124 42073 48127
rect 42024 48096 42073 48124
rect 42024 48084 42030 48096
rect 42061 48093 42073 48096
rect 42107 48093 42119 48127
rect 42061 48087 42119 48093
rect 42245 48127 42303 48133
rect 42245 48093 42257 48127
rect 42291 48093 42303 48127
rect 42245 48087 42303 48093
rect 42705 48127 42763 48133
rect 42705 48093 42717 48127
rect 42751 48124 42763 48127
rect 43990 48124 43996 48136
rect 42751 48096 43996 48124
rect 42751 48093 42763 48096
rect 42705 48087 42763 48093
rect 43990 48084 43996 48096
rect 44048 48084 44054 48136
rect 45186 48124 45192 48136
rect 45147 48096 45192 48124
rect 45186 48084 45192 48096
rect 45244 48084 45250 48136
rect 45281 48127 45339 48133
rect 45281 48093 45293 48127
rect 45327 48093 45339 48127
rect 45281 48087 45339 48093
rect 40920 48028 41414 48056
rect 40920 48016 40926 48028
rect 42886 48016 42892 48068
rect 42944 48056 42950 48068
rect 44085 48059 44143 48065
rect 44085 48056 44097 48059
rect 42944 48028 44097 48056
rect 42944 48016 42950 48028
rect 44085 48025 44097 48028
rect 44131 48056 44143 48059
rect 45296 48056 45324 48087
rect 45370 48084 45376 48136
rect 45428 48124 45434 48136
rect 45480 48124 45508 48155
rect 46566 48152 46572 48204
rect 46624 48192 46630 48204
rect 56336 48201 56364 48232
rect 57238 48220 57244 48232
rect 57296 48220 57302 48272
rect 46937 48195 46995 48201
rect 46937 48192 46949 48195
rect 46624 48164 46949 48192
rect 46624 48152 46630 48164
rect 46937 48161 46949 48164
rect 46983 48161 46995 48195
rect 46937 48155 46995 48161
rect 56321 48195 56379 48201
rect 56321 48161 56333 48195
rect 56367 48161 56379 48195
rect 56321 48155 56379 48161
rect 56505 48195 56563 48201
rect 56505 48161 56517 48195
rect 56551 48192 56563 48195
rect 57146 48192 57152 48204
rect 56551 48164 57152 48192
rect 56551 48161 56563 48164
rect 56505 48155 56563 48161
rect 57146 48152 57152 48164
rect 57204 48152 57210 48204
rect 57882 48192 57888 48204
rect 57843 48164 57888 48192
rect 57882 48152 57888 48164
rect 57940 48152 57946 48204
rect 45428 48096 45508 48124
rect 45557 48127 45615 48133
rect 45428 48084 45434 48096
rect 45557 48093 45569 48127
rect 45603 48124 45615 48127
rect 46290 48124 46296 48136
rect 45603 48096 46152 48124
rect 46251 48096 46296 48124
rect 45603 48093 45615 48096
rect 45557 48087 45615 48093
rect 44131 48028 45324 48056
rect 44131 48025 44143 48028
rect 44085 48019 44143 48025
rect 45830 48016 45836 48068
rect 45888 48056 45894 48068
rect 46017 48059 46075 48065
rect 46017 48056 46029 48059
rect 45888 48028 46029 48056
rect 45888 48016 45894 48028
rect 46017 48025 46029 48028
rect 46063 48025 46075 48059
rect 46124 48056 46152 48096
rect 46290 48084 46296 48096
rect 46348 48084 46354 48136
rect 47029 48127 47087 48133
rect 47029 48093 47041 48127
rect 47075 48093 47087 48127
rect 47029 48087 47087 48093
rect 46382 48056 46388 48068
rect 46124 48028 46388 48056
rect 46017 48019 46075 48025
rect 46382 48016 46388 48028
rect 46440 48016 46446 48068
rect 46934 48016 46940 48068
rect 46992 48056 46998 48068
rect 47044 48056 47072 48087
rect 47394 48084 47400 48136
rect 47452 48124 47458 48136
rect 47949 48127 48007 48133
rect 47949 48124 47961 48127
rect 47452 48096 47961 48124
rect 47452 48084 47458 48096
rect 47949 48093 47961 48096
rect 47995 48093 48007 48127
rect 47949 48087 48007 48093
rect 48133 48127 48191 48133
rect 48133 48093 48145 48127
rect 48179 48093 48191 48127
rect 48133 48087 48191 48093
rect 46992 48028 47072 48056
rect 46992 48016 46998 48028
rect 47670 48016 47676 48068
rect 47728 48056 47734 48068
rect 48148 48056 48176 48087
rect 47728 48028 48176 48056
rect 47728 48016 47734 48028
rect 37424 47960 37964 47988
rect 37424 47948 37430 47960
rect 43622 47948 43628 48000
rect 43680 47988 43686 48000
rect 44177 47991 44235 47997
rect 44177 47988 44189 47991
rect 43680 47960 44189 47988
rect 43680 47948 43686 47960
rect 44177 47957 44189 47960
rect 44223 47957 44235 47991
rect 44177 47951 44235 47957
rect 45005 47991 45063 47997
rect 45005 47957 45017 47991
rect 45051 47988 45063 47991
rect 45462 47988 45468 48000
rect 45051 47960 45468 47988
rect 45051 47957 45063 47960
rect 45005 47951 45063 47957
rect 45462 47948 45468 47960
rect 45520 47948 45526 48000
rect 46198 47988 46204 48000
rect 46159 47960 46204 47988
rect 46198 47948 46204 47960
rect 46256 47948 46262 48000
rect 47397 47991 47455 47997
rect 47397 47957 47409 47991
rect 47443 47988 47455 47991
rect 47762 47988 47768 48000
rect 47443 47960 47768 47988
rect 47443 47957 47455 47960
rect 47397 47951 47455 47957
rect 47762 47948 47768 47960
rect 47820 47948 47826 48000
rect 48133 47991 48191 47997
rect 48133 47957 48145 47991
rect 48179 47988 48191 47991
rect 48774 47988 48780 48000
rect 48179 47960 48780 47988
rect 48179 47957 48191 47960
rect 48133 47951 48191 47957
rect 48774 47948 48780 47960
rect 48832 47948 48838 48000
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 20625 47787 20683 47793
rect 20625 47753 20637 47787
rect 20671 47753 20683 47787
rect 24670 47784 24676 47796
rect 20625 47747 20683 47753
rect 24320 47756 24676 47784
rect 19052 47719 19110 47725
rect 19052 47685 19064 47719
rect 19098 47716 19110 47719
rect 20640 47716 20668 47747
rect 24320 47725 24348 47756
rect 24670 47744 24676 47756
rect 24728 47744 24734 47796
rect 33042 47784 33048 47796
rect 33003 47756 33048 47784
rect 33042 47744 33048 47756
rect 33100 47744 33106 47796
rect 33870 47744 33876 47796
rect 33928 47784 33934 47796
rect 37826 47784 37832 47796
rect 33928 47756 37688 47784
rect 37787 47756 37832 47784
rect 33928 47744 33934 47756
rect 19098 47688 20668 47716
rect 24305 47719 24363 47725
rect 19098 47685 19110 47688
rect 19052 47679 19110 47685
rect 24305 47685 24317 47719
rect 24351 47685 24363 47719
rect 24305 47679 24363 47685
rect 24535 47719 24593 47725
rect 24535 47685 24547 47719
rect 24581 47716 24593 47719
rect 24762 47716 24768 47728
rect 24581 47688 24768 47716
rect 24581 47685 24593 47688
rect 24535 47679 24593 47685
rect 24762 47676 24768 47688
rect 24820 47676 24826 47728
rect 25869 47719 25927 47725
rect 25869 47685 25881 47719
rect 25915 47716 25927 47719
rect 29546 47716 29552 47728
rect 25915 47688 29552 47716
rect 25915 47685 25927 47688
rect 25869 47679 25927 47685
rect 29546 47676 29552 47688
rect 29604 47716 29610 47728
rect 29733 47719 29791 47725
rect 29733 47716 29745 47719
rect 29604 47688 29745 47716
rect 29604 47676 29610 47688
rect 29733 47685 29745 47688
rect 29779 47685 29791 47719
rect 29733 47679 29791 47685
rect 29917 47719 29975 47725
rect 29917 47685 29929 47719
rect 29963 47716 29975 47719
rect 30558 47716 30564 47728
rect 29963 47688 30564 47716
rect 29963 47685 29975 47688
rect 29917 47679 29975 47685
rect 30558 47676 30564 47688
rect 30616 47676 30622 47728
rect 37550 47716 37556 47728
rect 30668 47688 35204 47716
rect 37511 47688 37556 47716
rect 8938 47608 8944 47660
rect 8996 47648 9002 47660
rect 20806 47648 20812 47660
rect 8996 47620 19840 47648
rect 20767 47620 20812 47648
rect 8996 47608 9002 47620
rect 18782 47580 18788 47592
rect 18743 47552 18788 47580
rect 18782 47540 18788 47552
rect 18840 47540 18846 47592
rect 19812 47580 19840 47620
rect 20806 47608 20812 47620
rect 20864 47608 20870 47660
rect 24210 47648 24216 47660
rect 24171 47620 24216 47648
rect 24210 47608 24216 47620
rect 24268 47608 24274 47660
rect 24397 47651 24455 47657
rect 24397 47617 24409 47651
rect 24443 47648 24455 47651
rect 26050 47648 26056 47660
rect 24443 47620 26056 47648
rect 24443 47617 24455 47620
rect 24397 47611 24455 47617
rect 26050 47608 26056 47620
rect 26108 47608 26114 47660
rect 26142 47608 26148 47660
rect 26200 47648 26206 47660
rect 27433 47651 27491 47657
rect 27433 47648 27445 47651
rect 26200 47620 27445 47648
rect 26200 47608 26206 47620
rect 27433 47617 27445 47620
rect 27479 47617 27491 47651
rect 27614 47648 27620 47660
rect 27575 47620 27620 47648
rect 27433 47611 27491 47617
rect 27614 47608 27620 47620
rect 27672 47608 27678 47660
rect 28258 47648 28264 47660
rect 28219 47620 28264 47648
rect 28258 47608 28264 47620
rect 28316 47608 28322 47660
rect 30374 47648 30380 47660
rect 30335 47620 30380 47648
rect 30374 47608 30380 47620
rect 30432 47648 30438 47660
rect 30668 47648 30696 47688
rect 30432 47620 30696 47648
rect 31113 47651 31171 47657
rect 30432 47608 30438 47620
rect 31113 47617 31125 47651
rect 31159 47617 31171 47651
rect 31113 47611 31171 47617
rect 24670 47580 24676 47592
rect 19812 47552 22094 47580
rect 24631 47552 24676 47580
rect 22066 47512 22094 47552
rect 24670 47540 24676 47552
rect 24728 47540 24734 47592
rect 28902 47580 28908 47592
rect 28863 47552 28908 47580
rect 28902 47540 28908 47552
rect 28960 47540 28966 47592
rect 30466 47540 30472 47592
rect 30524 47580 30530 47592
rect 31128 47580 31156 47611
rect 31938 47608 31944 47660
rect 31996 47648 32002 47660
rect 32309 47651 32367 47657
rect 32309 47648 32321 47651
rect 31996 47620 32321 47648
rect 31996 47608 32002 47620
rect 32309 47617 32321 47620
rect 32355 47617 32367 47651
rect 32309 47611 32367 47617
rect 32398 47608 32404 47660
rect 32456 47648 32462 47660
rect 32493 47651 32551 47657
rect 32493 47648 32505 47651
rect 32456 47620 32505 47648
rect 32456 47608 32462 47620
rect 32493 47617 32505 47620
rect 32539 47617 32551 47651
rect 32493 47611 32551 47617
rect 32508 47580 32536 47611
rect 32582 47608 32588 47660
rect 32640 47648 32646 47660
rect 33318 47648 33324 47660
rect 32640 47620 32685 47648
rect 33279 47620 33324 47648
rect 32640 47608 32646 47620
rect 33318 47608 33324 47620
rect 33376 47608 33382 47660
rect 33413 47651 33471 47657
rect 33413 47617 33425 47651
rect 33459 47617 33471 47651
rect 33413 47611 33471 47617
rect 33428 47580 33456 47611
rect 33502 47608 33508 47660
rect 33560 47648 33566 47660
rect 33686 47648 33692 47660
rect 33560 47620 33605 47648
rect 33647 47620 33692 47648
rect 33560 47608 33566 47620
rect 33686 47608 33692 47620
rect 33744 47608 33750 47660
rect 34146 47648 34152 47660
rect 34107 47620 34152 47648
rect 34146 47608 34152 47620
rect 34204 47608 34210 47660
rect 34405 47651 34463 47657
rect 34405 47648 34417 47651
rect 34256 47620 34417 47648
rect 34256 47580 34284 47620
rect 34405 47617 34417 47620
rect 34451 47617 34463 47651
rect 34405 47611 34463 47617
rect 30524 47552 32076 47580
rect 32508 47552 33456 47580
rect 34164 47552 34284 47580
rect 35176 47580 35204 47688
rect 37550 47676 37556 47688
rect 37608 47676 37614 47728
rect 37274 47648 37280 47660
rect 37235 47620 37280 47648
rect 37274 47608 37280 47620
rect 37332 47608 37338 47660
rect 37366 47608 37372 47660
rect 37424 47648 37430 47660
rect 37660 47657 37688 47756
rect 37826 47744 37832 47756
rect 37884 47744 37890 47796
rect 40037 47787 40095 47793
rect 40037 47753 40049 47787
rect 40083 47784 40095 47787
rect 44545 47787 44603 47793
rect 40083 47756 41460 47784
rect 40083 47753 40095 47756
rect 40037 47747 40095 47753
rect 40586 47716 40592 47728
rect 40547 47688 40592 47716
rect 40586 47676 40592 47688
rect 40644 47676 40650 47728
rect 41432 47660 41460 47756
rect 44545 47753 44557 47787
rect 44591 47784 44603 47787
rect 44910 47784 44916 47796
rect 44591 47756 44916 47784
rect 44591 47753 44603 47756
rect 44545 47747 44603 47753
rect 44910 47744 44916 47756
rect 44968 47744 44974 47796
rect 45186 47744 45192 47796
rect 45244 47784 45250 47796
rect 46106 47784 46112 47796
rect 45244 47756 46112 47784
rect 45244 47744 45250 47756
rect 46106 47744 46112 47756
rect 46164 47744 46170 47796
rect 46477 47787 46535 47793
rect 46477 47753 46489 47787
rect 46523 47784 46535 47787
rect 46934 47784 46940 47796
rect 46523 47756 46940 47784
rect 46523 47753 46535 47756
rect 46477 47747 46535 47753
rect 46934 47744 46940 47756
rect 46992 47744 46998 47796
rect 44082 47676 44088 47728
rect 44140 47716 44146 47728
rect 45005 47719 45063 47725
rect 44140 47688 44496 47716
rect 44140 47676 44146 47688
rect 37461 47651 37519 47657
rect 37461 47648 37473 47651
rect 37424 47620 37473 47648
rect 37424 47608 37430 47620
rect 37461 47617 37473 47620
rect 37507 47617 37519 47651
rect 37461 47611 37519 47617
rect 37645 47651 37703 47657
rect 37645 47617 37657 47651
rect 37691 47648 37703 47651
rect 38102 47648 38108 47660
rect 37691 47620 38108 47648
rect 37691 47617 37703 47620
rect 37645 47611 37703 47617
rect 38102 47608 38108 47620
rect 38160 47608 38166 47660
rect 39206 47608 39212 47660
rect 39264 47648 39270 47660
rect 39577 47651 39635 47657
rect 39577 47648 39589 47651
rect 39264 47620 39589 47648
rect 39264 47608 39270 47620
rect 39577 47617 39589 47620
rect 39623 47617 39635 47651
rect 39577 47611 39635 47617
rect 41138 47608 41144 47660
rect 41196 47648 41202 47660
rect 41325 47651 41383 47657
rect 41325 47648 41337 47651
rect 41196 47620 41337 47648
rect 41196 47608 41202 47620
rect 41325 47617 41337 47620
rect 41371 47617 41383 47651
rect 41325 47611 41383 47617
rect 41414 47608 41420 47660
rect 41472 47648 41478 47660
rect 41509 47651 41567 47657
rect 41509 47648 41521 47651
rect 41472 47620 41521 47648
rect 41472 47608 41478 47620
rect 41509 47617 41521 47620
rect 41555 47617 41567 47651
rect 44174 47648 44180 47660
rect 44135 47620 44180 47648
rect 41509 47611 41567 47617
rect 44174 47608 44180 47620
rect 44232 47608 44238 47660
rect 44361 47651 44419 47657
rect 44361 47617 44373 47651
rect 44407 47617 44419 47651
rect 44468 47648 44496 47688
rect 45005 47685 45017 47719
rect 45051 47716 45063 47719
rect 45051 47688 48084 47716
rect 45051 47685 45063 47688
rect 45005 47679 45063 47685
rect 44910 47648 44916 47660
rect 44468 47620 44916 47648
rect 44361 47611 44419 47617
rect 44266 47580 44272 47592
rect 35176 47552 44272 47580
rect 30524 47540 30530 47552
rect 28920 47512 28948 47540
rect 22066 47484 28948 47512
rect 19518 47404 19524 47456
rect 19576 47444 19582 47456
rect 20162 47444 20168 47456
rect 19576 47416 20168 47444
rect 19576 47404 19582 47416
rect 20162 47404 20168 47416
rect 20220 47404 20226 47456
rect 24029 47447 24087 47453
rect 24029 47413 24041 47447
rect 24075 47444 24087 47447
rect 24486 47444 24492 47456
rect 24075 47416 24492 47444
rect 24075 47413 24087 47416
rect 24029 47407 24087 47413
rect 24486 47404 24492 47416
rect 24544 47404 24550 47456
rect 25958 47444 25964 47456
rect 25919 47416 25964 47444
rect 25958 47404 25964 47416
rect 26016 47404 26022 47456
rect 27614 47404 27620 47456
rect 27672 47444 27678 47456
rect 30469 47447 30527 47453
rect 30469 47444 30481 47447
rect 27672 47416 30481 47444
rect 27672 47404 27678 47416
rect 30469 47413 30481 47416
rect 30515 47413 30527 47447
rect 30469 47407 30527 47413
rect 31205 47447 31263 47453
rect 31205 47413 31217 47447
rect 31251 47444 31263 47447
rect 31846 47444 31852 47456
rect 31251 47416 31852 47444
rect 31251 47413 31263 47416
rect 31205 47407 31263 47413
rect 31846 47404 31852 47416
rect 31904 47404 31910 47456
rect 32048 47444 32076 47552
rect 32125 47515 32183 47521
rect 32125 47481 32137 47515
rect 32171 47512 32183 47515
rect 34164 47512 34192 47552
rect 44266 47540 44272 47552
rect 44324 47540 44330 47592
rect 44376 47580 44404 47611
rect 44910 47608 44916 47620
rect 44968 47648 44974 47660
rect 45235 47651 45293 47657
rect 45235 47648 45247 47651
rect 44968 47620 45247 47648
rect 44968 47608 44974 47620
rect 45235 47617 45247 47620
rect 45281 47617 45293 47651
rect 45370 47648 45376 47660
rect 45331 47620 45376 47648
rect 45235 47611 45293 47617
rect 45370 47608 45376 47620
rect 45428 47608 45434 47660
rect 45462 47608 45468 47660
rect 45520 47648 45526 47660
rect 45646 47648 45652 47660
rect 45520 47620 45565 47648
rect 45607 47620 45652 47648
rect 45520 47608 45526 47620
rect 45646 47608 45652 47620
rect 45704 47608 45710 47660
rect 46198 47648 46204 47660
rect 45756 47620 46204 47648
rect 45756 47580 45784 47620
rect 46198 47608 46204 47620
rect 46256 47608 46262 47660
rect 46566 47648 46572 47660
rect 46527 47620 46572 47648
rect 46566 47608 46572 47620
rect 46624 47608 46630 47660
rect 47854 47648 47860 47660
rect 47815 47620 47860 47648
rect 47854 47608 47860 47620
rect 47912 47608 47918 47660
rect 48056 47657 48084 47688
rect 47946 47651 48004 47657
rect 47946 47617 47958 47651
rect 47992 47617 48004 47651
rect 47946 47611 48004 47617
rect 48041 47651 48099 47657
rect 48041 47617 48053 47651
rect 48087 47617 48099 47651
rect 48222 47648 48228 47660
rect 48183 47620 48228 47648
rect 48041 47611 48099 47617
rect 46106 47580 46112 47592
rect 44376 47552 45784 47580
rect 46019 47552 46112 47580
rect 46106 47540 46112 47552
rect 46164 47580 46170 47592
rect 47026 47580 47032 47592
rect 46164 47552 47032 47580
rect 46164 47540 46170 47552
rect 47026 47540 47032 47552
rect 47084 47540 47090 47592
rect 47762 47540 47768 47592
rect 47820 47580 47826 47592
rect 47961 47580 47989 47611
rect 48222 47608 48228 47620
rect 48280 47608 48286 47660
rect 48406 47608 48412 47660
rect 48464 47648 48470 47660
rect 48869 47651 48927 47657
rect 48869 47648 48881 47651
rect 48464 47620 48881 47648
rect 48464 47608 48470 47620
rect 48869 47617 48881 47620
rect 48915 47617 48927 47651
rect 48869 47611 48927 47617
rect 48774 47580 48780 47592
rect 47820 47552 47989 47580
rect 48735 47552 48780 47580
rect 47820 47540 47826 47552
rect 48774 47540 48780 47552
rect 48832 47540 48838 47592
rect 35434 47512 35440 47524
rect 32171 47484 34192 47512
rect 35360 47484 35440 47512
rect 32171 47481 32183 47484
rect 32125 47475 32183 47481
rect 35360 47444 35388 47484
rect 35434 47472 35440 47484
rect 35492 47472 35498 47524
rect 39850 47512 39856 47524
rect 39811 47484 39856 47512
rect 39850 47472 39856 47484
rect 39908 47472 39914 47524
rect 44174 47472 44180 47524
rect 44232 47512 44238 47524
rect 46290 47512 46296 47524
rect 44232 47484 46296 47512
rect 44232 47472 44238 47484
rect 46290 47472 46296 47484
rect 46348 47472 46354 47524
rect 35526 47444 35532 47456
rect 32048 47416 35388 47444
rect 35487 47416 35532 47444
rect 35526 47404 35532 47416
rect 35584 47404 35590 47456
rect 37550 47404 37556 47456
rect 37608 47444 37614 47456
rect 40681 47447 40739 47453
rect 40681 47444 40693 47447
rect 37608 47416 40693 47444
rect 37608 47404 37614 47416
rect 40681 47413 40693 47416
rect 40727 47444 40739 47447
rect 40862 47444 40868 47456
rect 40727 47416 40868 47444
rect 40727 47413 40739 47416
rect 40681 47407 40739 47413
rect 40862 47404 40868 47416
rect 40920 47404 40926 47456
rect 41690 47444 41696 47456
rect 41603 47416 41696 47444
rect 41690 47404 41696 47416
rect 41748 47444 41754 47456
rect 45922 47444 45928 47456
rect 41748 47416 45928 47444
rect 41748 47404 41754 47416
rect 45922 47404 45928 47416
rect 45980 47404 45986 47456
rect 46106 47404 46112 47456
rect 46164 47444 46170 47456
rect 46566 47444 46572 47456
rect 46164 47416 46572 47444
rect 46164 47404 46170 47416
rect 46566 47404 46572 47416
rect 46624 47404 46630 47456
rect 47581 47447 47639 47453
rect 47581 47413 47593 47447
rect 47627 47444 47639 47447
rect 48774 47444 48780 47456
rect 47627 47416 48780 47444
rect 47627 47413 47639 47416
rect 47581 47407 47639 47413
rect 48774 47404 48780 47416
rect 48832 47404 48838 47456
rect 48866 47404 48872 47456
rect 48924 47444 48930 47456
rect 49145 47447 49203 47453
rect 49145 47444 49157 47447
rect 48924 47416 49157 47444
rect 48924 47404 48930 47416
rect 49145 47413 49157 47416
rect 49191 47413 49203 47447
rect 49145 47407 49203 47413
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 2958 47200 2964 47252
rect 3016 47240 3022 47252
rect 40954 47240 40960 47252
rect 3016 47212 27752 47240
rect 3016 47200 3022 47212
rect 19518 47104 19524 47116
rect 19479 47076 19524 47104
rect 19518 47064 19524 47076
rect 19576 47064 19582 47116
rect 20070 47064 20076 47116
rect 20128 47104 20134 47116
rect 20717 47107 20775 47113
rect 20717 47104 20729 47107
rect 20128 47076 20729 47104
rect 20128 47064 20134 47076
rect 20717 47073 20729 47076
rect 20763 47073 20775 47107
rect 27341 47107 27399 47113
rect 20717 47067 20775 47073
rect 20824 47076 24256 47104
rect 19334 46996 19340 47048
rect 19392 47036 19398 47048
rect 19705 47039 19763 47045
rect 19705 47036 19717 47039
rect 19392 47008 19717 47036
rect 19392 46996 19398 47008
rect 19705 47005 19717 47008
rect 19751 47036 19763 47039
rect 19978 47036 19984 47048
rect 19751 47008 19984 47036
rect 19751 47005 19763 47008
rect 19705 46999 19763 47005
rect 19978 46996 19984 47008
rect 20036 47036 20042 47048
rect 20346 47036 20352 47048
rect 20036 47008 20208 47036
rect 20307 47008 20352 47036
rect 20036 46996 20042 47008
rect 19426 46928 19432 46980
rect 19484 46968 19490 46980
rect 19889 46971 19947 46977
rect 19889 46968 19901 46971
rect 19484 46940 19901 46968
rect 19484 46928 19490 46940
rect 19889 46937 19901 46940
rect 19935 46937 19947 46971
rect 20180 46968 20208 47008
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 20533 47039 20591 47045
rect 20533 47005 20545 47039
rect 20579 47036 20591 47039
rect 20824 47036 20852 47076
rect 21358 47036 21364 47048
rect 20579 47008 20852 47036
rect 21319 47008 21364 47036
rect 20579 47005 20591 47008
rect 20533 46999 20591 47005
rect 20548 46968 20576 46999
rect 21358 46996 21364 47008
rect 21416 46996 21422 47048
rect 22833 47039 22891 47045
rect 22833 47005 22845 47039
rect 22879 47036 22891 47039
rect 24026 47036 24032 47048
rect 22879 47008 24032 47036
rect 22879 47005 22891 47008
rect 22833 46999 22891 47005
rect 24026 46996 24032 47008
rect 24084 46996 24090 47048
rect 20180 46940 20576 46968
rect 19889 46931 19947 46937
rect 20622 46928 20628 46980
rect 20680 46968 20686 46980
rect 21177 46971 21235 46977
rect 21177 46968 21189 46971
rect 20680 46940 21189 46968
rect 20680 46928 20686 46940
rect 21177 46937 21189 46940
rect 21223 46937 21235 46971
rect 21177 46931 21235 46937
rect 21545 46971 21603 46977
rect 21545 46937 21557 46971
rect 21591 46968 21603 46971
rect 22278 46968 22284 46980
rect 21591 46940 22284 46968
rect 21591 46937 21603 46940
rect 21545 46931 21603 46937
rect 22278 46928 22284 46940
rect 22336 46928 22342 46980
rect 24228 46968 24256 47076
rect 27341 47073 27353 47107
rect 27387 47104 27399 47107
rect 27614 47104 27620 47116
rect 27387 47076 27620 47104
rect 27387 47073 27399 47076
rect 27341 47067 27399 47073
rect 27614 47064 27620 47076
rect 27672 47064 27678 47116
rect 27724 47113 27752 47212
rect 35084 47212 40960 47240
rect 35084 47184 35112 47212
rect 40954 47200 40960 47212
rect 41012 47200 41018 47252
rect 41322 47200 41328 47252
rect 41380 47240 41386 47252
rect 41380 47212 41736 47240
rect 41380 47200 41386 47212
rect 30006 47172 30012 47184
rect 29967 47144 30012 47172
rect 30006 47132 30012 47144
rect 30064 47172 30070 47184
rect 30282 47172 30288 47184
rect 30064 47144 30288 47172
rect 30064 47132 30070 47144
rect 30282 47132 30288 47144
rect 30340 47132 30346 47184
rect 31018 47172 31024 47184
rect 30979 47144 31024 47172
rect 31018 47132 31024 47144
rect 31076 47132 31082 47184
rect 35066 47132 35072 47184
rect 35124 47132 35130 47184
rect 37274 47132 37280 47184
rect 37332 47172 37338 47184
rect 37642 47172 37648 47184
rect 37332 47144 37648 47172
rect 37332 47132 37338 47144
rect 37642 47132 37648 47144
rect 37700 47132 37706 47184
rect 39758 47132 39764 47184
rect 39816 47172 39822 47184
rect 41708 47172 41736 47212
rect 45370 47200 45376 47252
rect 45428 47240 45434 47252
rect 46017 47243 46075 47249
rect 46017 47240 46029 47243
rect 45428 47212 46029 47240
rect 45428 47200 45434 47212
rect 46017 47209 46029 47212
rect 46063 47209 46075 47243
rect 47946 47240 47952 47252
rect 47907 47212 47952 47240
rect 46017 47203 46075 47209
rect 47946 47200 47952 47212
rect 48004 47200 48010 47252
rect 48222 47240 48228 47252
rect 48183 47212 48228 47240
rect 48222 47200 48228 47212
rect 48280 47200 48286 47252
rect 56226 47172 56232 47184
rect 39816 47144 41644 47172
rect 41708 47144 56232 47172
rect 39816 47132 39822 47144
rect 27709 47107 27767 47113
rect 27709 47073 27721 47107
rect 27755 47073 27767 47107
rect 30098 47104 30104 47116
rect 30059 47076 30104 47104
rect 27709 47067 27767 47073
rect 30098 47064 30104 47076
rect 30156 47064 30162 47116
rect 30650 47064 30656 47116
rect 30708 47104 30714 47116
rect 31665 47107 31723 47113
rect 31665 47104 31677 47107
rect 30708 47076 31677 47104
rect 30708 47064 30714 47076
rect 31665 47073 31677 47076
rect 31711 47073 31723 47107
rect 31846 47104 31852 47116
rect 31807 47076 31852 47104
rect 31665 47067 31723 47073
rect 31846 47064 31852 47076
rect 31904 47064 31910 47116
rect 33502 47104 33508 47116
rect 33463 47076 33508 47104
rect 33502 47064 33508 47076
rect 33560 47064 33566 47116
rect 35434 47064 35440 47116
rect 35492 47104 35498 47116
rect 41322 47104 41328 47116
rect 35492 47076 41328 47104
rect 35492 47064 35498 47076
rect 41322 47064 41328 47076
rect 41380 47064 41386 47116
rect 24394 47036 24400 47048
rect 24355 47008 24400 47036
rect 24394 46996 24400 47008
rect 24452 46996 24458 47048
rect 24486 46996 24492 47048
rect 24544 47036 24550 47048
rect 24653 47039 24711 47045
rect 24653 47036 24665 47039
rect 24544 47008 24665 47036
rect 24544 46996 24550 47008
rect 24653 47005 24665 47008
rect 24699 47005 24711 47039
rect 24653 46999 24711 47005
rect 26142 46996 26148 47048
rect 26200 47036 26206 47048
rect 26237 47039 26295 47045
rect 26237 47036 26249 47039
rect 26200 47008 26249 47036
rect 26200 46996 26206 47008
rect 26237 47005 26249 47008
rect 26283 47005 26295 47039
rect 27154 47036 27160 47048
rect 27115 47008 27160 47036
rect 26237 46999 26295 47005
rect 27154 46996 27160 47008
rect 27212 46996 27218 47048
rect 30558 46996 30564 47048
rect 30616 47036 30622 47048
rect 30837 47039 30895 47045
rect 30837 47036 30849 47039
rect 30616 47008 30849 47036
rect 30616 46996 30622 47008
rect 30837 47005 30849 47008
rect 30883 47005 30895 47039
rect 35066 47036 35072 47048
rect 35027 47008 35072 47036
rect 30837 46999 30895 47005
rect 35066 46996 35072 47008
rect 35124 46996 35130 47048
rect 35253 47039 35311 47045
rect 35253 47005 35265 47039
rect 35299 47005 35311 47039
rect 35253 46999 35311 47005
rect 27614 46968 27620 46980
rect 24228 46940 27620 46968
rect 27614 46928 27620 46940
rect 27672 46928 27678 46980
rect 29641 46971 29699 46977
rect 29641 46937 29653 46971
rect 29687 46968 29699 46971
rect 31386 46968 31392 46980
rect 29687 46940 31392 46968
rect 29687 46937 29699 46940
rect 29641 46931 29699 46937
rect 31386 46928 31392 46940
rect 31444 46928 31450 46980
rect 33594 46928 33600 46980
rect 33652 46968 33658 46980
rect 35161 46971 35219 46977
rect 35161 46968 35173 46971
rect 33652 46940 35173 46968
rect 33652 46928 33658 46940
rect 35161 46937 35173 46940
rect 35207 46937 35219 46971
rect 35161 46931 35219 46937
rect 22646 46900 22652 46912
rect 22607 46872 22652 46900
rect 22646 46860 22652 46872
rect 22704 46860 22710 46912
rect 25774 46900 25780 46912
rect 25735 46872 25780 46900
rect 25774 46860 25780 46872
rect 25832 46860 25838 46912
rect 26421 46903 26479 46909
rect 26421 46869 26433 46903
rect 26467 46900 26479 46903
rect 26970 46900 26976 46912
rect 26467 46872 26976 46900
rect 26467 46869 26479 46872
rect 26421 46863 26479 46869
rect 26970 46860 26976 46872
rect 27028 46860 27034 46912
rect 34698 46860 34704 46912
rect 34756 46900 34762 46912
rect 35268 46900 35296 46999
rect 35894 46996 35900 47048
rect 35952 47036 35958 47048
rect 36449 47039 36507 47045
rect 36449 47036 36461 47039
rect 35952 47008 36461 47036
rect 35952 46996 35958 47008
rect 36449 47005 36461 47008
rect 36495 47005 36507 47039
rect 39666 47036 39672 47048
rect 36449 46999 36507 47005
rect 37844 47008 39672 47036
rect 35526 46928 35532 46980
rect 35584 46968 35590 46980
rect 36265 46971 36323 46977
rect 36265 46968 36277 46971
rect 35584 46940 36277 46968
rect 35584 46928 35590 46940
rect 36265 46937 36277 46940
rect 36311 46968 36323 46971
rect 37844 46968 37872 47008
rect 39666 46996 39672 47008
rect 39724 46996 39730 47048
rect 39758 46996 39764 47048
rect 39816 47036 39822 47048
rect 39945 47039 40003 47045
rect 39945 47036 39957 47039
rect 39816 47008 39957 47036
rect 39816 46996 39822 47008
rect 39945 47005 39957 47008
rect 39991 47005 40003 47039
rect 39945 46999 40003 47005
rect 40037 47039 40095 47045
rect 40037 47005 40049 47039
rect 40083 47005 40095 47039
rect 40037 46999 40095 47005
rect 40221 47039 40279 47045
rect 40221 47005 40233 47039
rect 40267 47005 40279 47039
rect 40221 46999 40279 47005
rect 36311 46940 37872 46968
rect 36311 46937 36323 46940
rect 36265 46931 36323 46937
rect 37918 46928 37924 46980
rect 37976 46968 37982 46980
rect 40052 46968 40080 46999
rect 37976 46940 40080 46968
rect 40236 46968 40264 46999
rect 40310 46996 40316 47048
rect 40368 47036 40374 47048
rect 41414 47036 41420 47048
rect 40368 47008 40413 47036
rect 40368 46996 40374 47008
rect 41386 46996 41420 47036
rect 41472 47036 41478 47048
rect 41616 47045 41644 47144
rect 56226 47132 56232 47144
rect 56284 47132 56290 47184
rect 44910 47064 44916 47116
rect 44968 47104 44974 47116
rect 46753 47107 46811 47113
rect 44968 47076 45600 47104
rect 44968 47064 44974 47076
rect 41601 47039 41659 47045
rect 41472 47008 41517 47036
rect 41472 46996 41478 47008
rect 41601 47005 41613 47039
rect 41647 47036 41659 47039
rect 42337 47039 42395 47045
rect 42337 47036 42349 47039
rect 41647 47008 42349 47036
rect 41647 47005 41659 47008
rect 41601 46999 41659 47005
rect 42337 47005 42349 47008
rect 42383 47005 42395 47039
rect 42337 46999 42395 47005
rect 42886 46996 42892 47048
rect 42944 47036 42950 47048
rect 44453 47039 44511 47045
rect 44453 47036 44465 47039
rect 42944 47008 44465 47036
rect 42944 46996 42950 47008
rect 44453 47005 44465 47008
rect 44499 47005 44511 47039
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 44453 46999 44511 47005
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 45281 47039 45339 47045
rect 45281 47005 45293 47039
rect 45327 47036 45339 47039
rect 45370 47036 45376 47048
rect 45327 47008 45376 47036
rect 45327 47005 45339 47008
rect 45281 46999 45339 47005
rect 45370 46996 45376 47008
rect 45428 46996 45434 47048
rect 45572 47045 45600 47076
rect 46753 47073 46765 47107
rect 46799 47104 46811 47107
rect 49145 47107 49203 47113
rect 46799 47076 47716 47104
rect 46799 47073 46811 47076
rect 46753 47067 46811 47073
rect 47688 47048 47716 47076
rect 48286 47076 49004 47104
rect 45465 47039 45523 47045
rect 45465 47005 45477 47039
rect 45511 47005 45523 47039
rect 45465 46999 45523 47005
rect 45557 47039 45615 47045
rect 45557 47005 45569 47039
rect 45603 47005 45615 47039
rect 45557 46999 45615 47005
rect 41386 46968 41414 46996
rect 40236 46940 41414 46968
rect 41693 46971 41751 46977
rect 37976 46928 37982 46940
rect 41693 46937 41705 46971
rect 41739 46968 41751 46971
rect 41966 46968 41972 46980
rect 41739 46940 41972 46968
rect 41739 46937 41751 46940
rect 41693 46931 41751 46937
rect 41966 46928 41972 46940
rect 42024 46928 42030 46980
rect 42153 46971 42211 46977
rect 42153 46937 42165 46971
rect 42199 46968 42211 46971
rect 42426 46968 42432 46980
rect 42199 46940 42432 46968
rect 42199 46937 42211 46940
rect 42153 46931 42211 46937
rect 40310 46900 40316 46912
rect 34756 46872 35296 46900
rect 40271 46872 40316 46900
rect 34756 46860 34762 46872
rect 40310 46860 40316 46872
rect 40368 46860 40374 46912
rect 41506 46860 41512 46912
rect 41564 46900 41570 46912
rect 42168 46900 42196 46931
rect 42426 46928 42432 46940
rect 42484 46928 42490 46980
rect 42521 46971 42579 46977
rect 42521 46937 42533 46971
rect 42567 46968 42579 46971
rect 42794 46968 42800 46980
rect 42567 46940 42800 46968
rect 42567 46937 42579 46940
rect 42521 46931 42579 46937
rect 42794 46928 42800 46940
rect 42852 46968 42858 46980
rect 43073 46971 43131 46977
rect 43073 46968 43085 46971
rect 42852 46940 43085 46968
rect 42852 46928 42858 46940
rect 43073 46937 43085 46940
rect 43119 46937 43131 46971
rect 43073 46931 43131 46937
rect 44085 46971 44143 46977
rect 44085 46937 44097 46971
rect 44131 46968 44143 46971
rect 44174 46968 44180 46980
rect 44131 46940 44180 46968
rect 44131 46937 44143 46940
rect 44085 46931 44143 46937
rect 44174 46928 44180 46940
rect 44232 46928 44238 46980
rect 44269 46971 44327 46977
rect 44269 46937 44281 46971
rect 44315 46968 44327 46971
rect 45480 46968 45508 46999
rect 45922 46996 45928 47048
rect 45980 47036 45986 47048
rect 46293 47039 46351 47045
rect 46293 47036 46305 47039
rect 45980 47008 46305 47036
rect 45980 46996 45986 47008
rect 46293 47005 46305 47008
rect 46339 47005 46351 47039
rect 46934 47036 46940 47048
rect 46847 47008 46940 47036
rect 46293 46999 46351 47005
rect 46934 46996 46940 47008
rect 46992 46996 46998 47048
rect 47118 47036 47124 47048
rect 47079 47008 47124 47036
rect 47118 46996 47124 47008
rect 47176 46996 47182 47048
rect 47210 46996 47216 47048
rect 47268 47036 47274 47048
rect 47670 47036 47676 47048
rect 47268 47008 47313 47036
rect 47631 47008 47676 47036
rect 47268 46996 47274 47008
rect 47670 46996 47676 47008
rect 47728 46996 47734 47048
rect 47854 46996 47860 47048
rect 47912 47036 47918 47048
rect 47949 47039 48007 47045
rect 47949 47036 47961 47039
rect 47912 47008 47961 47036
rect 47912 46996 47918 47008
rect 47949 47005 47961 47008
rect 47995 47036 48007 47039
rect 48286 47036 48314 47076
rect 48866 47036 48872 47048
rect 47995 47008 48314 47036
rect 48827 47008 48872 47036
rect 47995 47005 48007 47008
rect 47949 46999 48007 47005
rect 48866 46996 48872 47008
rect 48924 46996 48930 47048
rect 48976 47045 49004 47076
rect 49145 47073 49157 47107
rect 49191 47104 49203 47107
rect 50157 47107 50215 47113
rect 50157 47104 50169 47107
rect 49191 47076 50169 47104
rect 49191 47073 49203 47076
rect 49145 47067 49203 47073
rect 50157 47073 50169 47076
rect 50203 47073 50215 47107
rect 50157 47067 50215 47073
rect 56321 47107 56379 47113
rect 56321 47073 56333 47107
rect 56367 47104 56379 47107
rect 58066 47104 58072 47116
rect 56367 47076 58072 47104
rect 56367 47073 56379 47076
rect 56321 47067 56379 47073
rect 58066 47064 58072 47076
rect 58124 47064 58130 47116
rect 48961 47039 49019 47045
rect 48961 47005 48973 47039
rect 49007 47005 49019 47039
rect 48961 46999 49019 47005
rect 49237 47039 49295 47045
rect 49237 47005 49249 47039
rect 49283 47036 49295 47039
rect 49878 47036 49884 47048
rect 49283 47008 49884 47036
rect 49283 47005 49295 47008
rect 49237 46999 49295 47005
rect 49878 46996 49884 47008
rect 49936 46996 49942 47048
rect 49970 46996 49976 47048
rect 50028 47036 50034 47048
rect 50341 47039 50399 47045
rect 50341 47036 50353 47039
rect 50028 47008 50353 47036
rect 50028 46996 50034 47008
rect 50341 47005 50353 47008
rect 50387 47005 50399 47039
rect 50341 46999 50399 47005
rect 50617 47039 50675 47045
rect 50617 47005 50629 47039
rect 50663 47005 50675 47039
rect 50617 46999 50675 47005
rect 45738 46968 45744 46980
rect 44315 46940 45744 46968
rect 44315 46937 44327 46940
rect 44269 46931 44327 46937
rect 45738 46928 45744 46940
rect 45796 46928 45802 46980
rect 46017 46971 46075 46977
rect 46017 46937 46029 46971
rect 46063 46968 46075 46971
rect 46952 46968 46980 46996
rect 47762 46968 47768 46980
rect 46063 46940 47768 46968
rect 46063 46937 46075 46940
rect 46017 46931 46075 46937
rect 47762 46928 47768 46940
rect 47820 46928 47826 46980
rect 48314 46968 48320 46980
rect 47872 46940 48320 46968
rect 43162 46900 43168 46912
rect 41564 46872 42196 46900
rect 43123 46872 43168 46900
rect 41564 46860 41570 46872
rect 43162 46860 43168 46872
rect 43220 46860 43226 46912
rect 44726 46860 44732 46912
rect 44784 46900 44790 46912
rect 45005 46903 45063 46909
rect 45005 46900 45017 46903
rect 44784 46872 45017 46900
rect 44784 46860 44790 46872
rect 45005 46869 45017 46872
rect 45051 46869 45063 46903
rect 45005 46863 45063 46869
rect 46201 46903 46259 46909
rect 46201 46869 46213 46903
rect 46247 46900 46259 46903
rect 46382 46900 46388 46912
rect 46247 46872 46388 46900
rect 46247 46869 46259 46872
rect 46201 46863 46259 46869
rect 46382 46860 46388 46872
rect 46440 46900 46446 46912
rect 47872 46900 47900 46940
rect 48314 46928 48320 46940
rect 48372 46928 48378 46980
rect 49786 46928 49792 46980
rect 49844 46968 49850 46980
rect 50632 46968 50660 46999
rect 49844 46940 50660 46968
rect 56505 46971 56563 46977
rect 49844 46928 49850 46940
rect 56505 46937 56517 46971
rect 56551 46968 56563 46971
rect 56962 46968 56968 46980
rect 56551 46940 56968 46968
rect 56551 46937 56563 46940
rect 56505 46931 56563 46937
rect 56962 46928 56968 46940
rect 57020 46928 57026 46980
rect 58158 46968 58164 46980
rect 58119 46940 58164 46968
rect 58158 46928 58164 46940
rect 58216 46928 58222 46980
rect 48682 46900 48688 46912
rect 46440 46872 47900 46900
rect 48643 46872 48688 46900
rect 46440 46860 46446 46872
rect 48682 46860 48688 46872
rect 48740 46860 48746 46912
rect 49602 46860 49608 46912
rect 49660 46900 49666 46912
rect 49970 46900 49976 46912
rect 49660 46872 49976 46900
rect 49660 46860 49666 46872
rect 49970 46860 49976 46872
rect 50028 46860 50034 46912
rect 50062 46860 50068 46912
rect 50120 46900 50126 46912
rect 50525 46903 50583 46909
rect 50525 46900 50537 46903
rect 50120 46872 50537 46900
rect 50120 46860 50126 46872
rect 50525 46869 50537 46872
rect 50571 46869 50583 46903
rect 50525 46863 50583 46869
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 24026 46696 24032 46708
rect 22204 46668 22784 46696
rect 23987 46668 24032 46696
rect 19328 46631 19386 46637
rect 19328 46597 19340 46631
rect 19374 46628 19386 46631
rect 19978 46628 19984 46640
rect 19374 46600 19984 46628
rect 19374 46597 19386 46600
rect 19328 46591 19386 46597
rect 19978 46588 19984 46600
rect 20036 46588 20042 46640
rect 22204 46637 22232 46668
rect 22189 46631 22247 46637
rect 22189 46597 22201 46631
rect 22235 46597 22247 46631
rect 22189 46591 22247 46597
rect 22278 46588 22284 46640
rect 22336 46637 22342 46640
rect 22336 46631 22365 46637
rect 22353 46597 22365 46631
rect 22336 46591 22365 46597
rect 22336 46588 22342 46591
rect 18782 46520 18788 46572
rect 18840 46560 18846 46572
rect 19061 46563 19119 46569
rect 19061 46560 19073 46563
rect 18840 46532 19073 46560
rect 18840 46520 18846 46532
rect 19061 46529 19073 46532
rect 19107 46529 19119 46563
rect 22002 46560 22008 46572
rect 21963 46532 22008 46560
rect 19061 46523 19119 46529
rect 22002 46520 22008 46532
rect 22060 46520 22066 46572
rect 22094 46520 22100 46572
rect 22152 46560 22158 46572
rect 22465 46563 22523 46569
rect 22152 46532 22197 46560
rect 22152 46520 22158 46532
rect 22465 46529 22477 46563
rect 22511 46560 22523 46563
rect 22646 46560 22652 46572
rect 22511 46532 22652 46560
rect 22511 46529 22523 46532
rect 22465 46523 22523 46529
rect 22646 46520 22652 46532
rect 22704 46520 22710 46572
rect 22756 46424 22784 46668
rect 24026 46656 24032 46668
rect 24084 46656 24090 46708
rect 24854 46656 24860 46708
rect 24912 46696 24918 46708
rect 25593 46699 25651 46705
rect 25593 46696 25605 46699
rect 24912 46668 25605 46696
rect 24912 46656 24918 46668
rect 25593 46665 25605 46668
rect 25639 46696 25651 46699
rect 26142 46696 26148 46708
rect 25639 46668 26148 46696
rect 25639 46665 25651 46668
rect 25593 46659 25651 46665
rect 26142 46656 26148 46668
rect 26200 46656 26206 46708
rect 27614 46696 27620 46708
rect 27575 46668 27620 46696
rect 27614 46656 27620 46668
rect 27672 46696 27678 46708
rect 30006 46696 30012 46708
rect 27672 46668 30012 46696
rect 27672 46656 27678 46668
rect 30006 46656 30012 46668
rect 30064 46656 30070 46708
rect 31386 46696 31392 46708
rect 31347 46668 31392 46696
rect 31386 46656 31392 46668
rect 31444 46656 31450 46708
rect 36170 46696 36176 46708
rect 31726 46668 36176 46696
rect 23017 46631 23075 46637
rect 23017 46597 23029 46631
rect 23063 46628 23075 46631
rect 25958 46628 25964 46640
rect 23063 46600 25964 46628
rect 23063 46597 23075 46600
rect 23017 46591 23075 46597
rect 25958 46588 25964 46600
rect 26016 46588 26022 46640
rect 26237 46631 26295 46637
rect 26237 46597 26249 46631
rect 26283 46628 26295 46631
rect 27525 46631 27583 46637
rect 27525 46628 27537 46631
rect 26283 46600 27537 46628
rect 26283 46597 26295 46600
rect 26237 46591 26295 46597
rect 27525 46597 27537 46600
rect 27571 46628 27583 46631
rect 27706 46628 27712 46640
rect 27571 46600 27712 46628
rect 27571 46597 27583 46600
rect 27525 46591 27583 46597
rect 27706 46588 27712 46600
rect 27764 46588 27770 46640
rect 31018 46628 31024 46640
rect 30024 46600 31024 46628
rect 23845 46563 23903 46569
rect 23845 46529 23857 46563
rect 23891 46560 23903 46563
rect 24765 46563 24823 46569
rect 24765 46560 24777 46563
rect 23891 46532 24777 46560
rect 23891 46529 23903 46532
rect 23845 46523 23903 46529
rect 24765 46529 24777 46532
rect 24811 46560 24823 46563
rect 24854 46560 24860 46572
rect 24811 46532 24860 46560
rect 24811 46529 24823 46532
rect 24765 46523 24823 46529
rect 24854 46520 24860 46532
rect 24912 46520 24918 46572
rect 25501 46563 25559 46569
rect 25501 46529 25513 46563
rect 25547 46560 25559 46563
rect 28258 46560 28264 46572
rect 25547 46532 26004 46560
rect 28219 46532 28264 46560
rect 25547 46529 25559 46532
rect 25501 46523 25559 46529
rect 25976 46504 26004 46532
rect 28258 46520 28264 46532
rect 28316 46520 28322 46572
rect 30024 46569 30052 46600
rect 31018 46588 31024 46600
rect 31076 46588 31082 46640
rect 30282 46569 30288 46572
rect 30009 46563 30067 46569
rect 30009 46529 30021 46563
rect 30055 46529 30067 46563
rect 30276 46560 30288 46569
rect 30243 46532 30288 46560
rect 30009 46523 30067 46529
rect 30276 46523 30288 46532
rect 30282 46520 30288 46523
rect 30340 46520 30346 46572
rect 23658 46492 23664 46504
rect 23619 46464 23664 46492
rect 23658 46452 23664 46464
rect 23716 46452 23722 46504
rect 24581 46495 24639 46501
rect 24581 46461 24593 46495
rect 24627 46492 24639 46495
rect 25130 46492 25136 46504
rect 24627 46464 25136 46492
rect 24627 46461 24639 46464
rect 24581 46455 24639 46461
rect 25130 46452 25136 46464
rect 25188 46492 25194 46504
rect 25774 46492 25780 46504
rect 25188 46464 25780 46492
rect 25188 46452 25194 46464
rect 25774 46452 25780 46464
rect 25832 46452 25838 46504
rect 25958 46452 25964 46504
rect 26016 46492 26022 46504
rect 27154 46492 27160 46504
rect 26016 46464 27160 46492
rect 26016 46452 26022 46464
rect 27154 46452 27160 46464
rect 27212 46452 27218 46504
rect 29365 46495 29423 46501
rect 29365 46461 29377 46495
rect 29411 46492 29423 46495
rect 29914 46492 29920 46504
rect 29411 46464 29920 46492
rect 29411 46461 29423 46464
rect 29365 46455 29423 46461
rect 29914 46452 29920 46464
rect 29972 46452 29978 46504
rect 26418 46424 26424 46436
rect 22756 46396 26424 46424
rect 26418 46384 26424 46396
rect 26476 46384 26482 46436
rect 20438 46356 20444 46368
rect 20399 46328 20444 46356
rect 20438 46316 20444 46328
rect 20496 46316 20502 46368
rect 21818 46356 21824 46368
rect 21779 46328 21824 46356
rect 21818 46316 21824 46328
rect 21876 46316 21882 46368
rect 23106 46356 23112 46368
rect 23067 46328 23112 46356
rect 23106 46316 23112 46328
rect 23164 46316 23170 46368
rect 24946 46356 24952 46368
rect 24907 46328 24952 46356
rect 24946 46316 24952 46328
rect 25004 46316 25010 46368
rect 29914 46316 29920 46368
rect 29972 46356 29978 46368
rect 31726 46356 31754 46668
rect 36170 46656 36176 46668
rect 36228 46656 36234 46708
rect 39298 46696 39304 46708
rect 39132 46668 39304 46696
rect 33410 46628 33416 46640
rect 32600 46600 33416 46628
rect 32600 46572 32628 46600
rect 33410 46588 33416 46600
rect 33468 46588 33474 46640
rect 35342 46588 35348 46640
rect 35400 46628 35406 46640
rect 39132 46628 39160 46668
rect 39298 46656 39304 46668
rect 39356 46656 39362 46708
rect 41046 46696 41052 46708
rect 40233 46668 41052 46696
rect 35400 46600 39160 46628
rect 35400 46588 35406 46600
rect 40233 46575 40261 46668
rect 41046 46656 41052 46668
rect 41104 46656 41110 46708
rect 42613 46699 42671 46705
rect 42613 46665 42625 46699
rect 42659 46696 42671 46699
rect 43346 46696 43352 46708
rect 42659 46668 43352 46696
rect 42659 46665 42671 46668
rect 42613 46659 42671 46665
rect 43346 46656 43352 46668
rect 43404 46656 43410 46708
rect 45094 46696 45100 46708
rect 45055 46668 45100 46696
rect 45094 46656 45100 46668
rect 45152 46656 45158 46708
rect 50062 46656 50068 46708
rect 50120 46696 50126 46708
rect 51077 46699 51135 46705
rect 51077 46696 51089 46699
rect 50120 46668 51089 46696
rect 50120 46656 50126 46668
rect 51077 46665 51089 46668
rect 51123 46665 51135 46699
rect 56962 46696 56968 46708
rect 56923 46668 56968 46696
rect 51077 46659 51135 46665
rect 56962 46656 56968 46668
rect 57020 46656 57026 46708
rect 42886 46628 42892 46640
rect 42720 46600 42892 46628
rect 32398 46560 32404 46572
rect 32311 46532 32404 46560
rect 32398 46520 32404 46532
rect 32456 46520 32462 46572
rect 32490 46563 32548 46569
rect 32490 46529 32502 46563
rect 32536 46529 32548 46563
rect 32490 46523 32548 46529
rect 32585 46566 32643 46572
rect 32585 46532 32597 46566
rect 32631 46532 32643 46566
rect 32585 46526 32643 46532
rect 32769 46563 32827 46569
rect 32769 46529 32781 46563
rect 32815 46560 32827 46563
rect 33594 46560 33600 46572
rect 32815 46532 33600 46560
rect 32815 46529 32827 46532
rect 32769 46523 32827 46529
rect 32416 46492 32444 46520
rect 32416 46464 32470 46492
rect 32122 46356 32128 46368
rect 29972 46328 31754 46356
rect 32083 46328 32128 46356
rect 29972 46316 29978 46328
rect 32122 46316 32128 46328
rect 32180 46316 32186 46368
rect 32442 46356 32470 46464
rect 32505 46424 32533 46523
rect 33594 46520 33600 46532
rect 33652 46520 33658 46572
rect 34149 46563 34207 46569
rect 34149 46529 34161 46563
rect 34195 46560 34207 46563
rect 34698 46560 34704 46572
rect 34195 46532 34704 46560
rect 34195 46529 34207 46532
rect 34149 46523 34207 46529
rect 34698 46520 34704 46532
rect 34756 46560 34762 46572
rect 36081 46563 36139 46569
rect 36081 46560 36093 46563
rect 34756 46532 36093 46560
rect 34756 46520 34762 46532
rect 36081 46529 36093 46532
rect 36127 46529 36139 46563
rect 36081 46523 36139 46529
rect 37274 46520 37280 46572
rect 37332 46560 37338 46572
rect 37918 46560 37924 46572
rect 37332 46532 37924 46560
rect 37332 46520 37338 46532
rect 37918 46520 37924 46532
rect 37976 46520 37982 46572
rect 38105 46563 38163 46569
rect 38105 46529 38117 46563
rect 38151 46529 38163 46563
rect 39206 46560 39212 46572
rect 39167 46532 39212 46560
rect 38105 46523 38163 46529
rect 34425 46495 34483 46501
rect 34425 46461 34437 46495
rect 34471 46461 34483 46495
rect 34425 46455 34483 46461
rect 35805 46495 35863 46501
rect 35805 46461 35817 46495
rect 35851 46492 35863 46495
rect 35894 46492 35900 46504
rect 35851 46464 35900 46492
rect 35851 46461 35863 46464
rect 35805 46455 35863 46461
rect 32582 46424 32588 46436
rect 32505 46396 32588 46424
rect 32582 46384 32588 46396
rect 32640 46384 32646 46436
rect 34440 46356 34468 46455
rect 35894 46452 35900 46464
rect 35952 46452 35958 46504
rect 38120 46492 38148 46523
rect 39206 46520 39212 46532
rect 39264 46520 39270 46572
rect 39393 46563 39451 46569
rect 39393 46529 39405 46563
rect 39439 46560 39451 46563
rect 39758 46560 39764 46572
rect 39439 46532 39764 46560
rect 39439 46529 39451 46532
rect 39393 46523 39451 46529
rect 39758 46520 39764 46532
rect 39816 46520 39822 46572
rect 40126 46560 40132 46572
rect 40087 46532 40132 46560
rect 40126 46520 40132 46532
rect 40184 46520 40190 46572
rect 40218 46569 40276 46575
rect 40218 46535 40230 46569
rect 40264 46535 40276 46569
rect 40218 46529 40276 46535
rect 40310 46520 40316 46572
rect 40368 46560 40374 46572
rect 40497 46563 40555 46569
rect 40368 46532 40413 46560
rect 40368 46520 40374 46532
rect 40497 46529 40509 46563
rect 40543 46560 40555 46563
rect 40862 46560 40868 46572
rect 40543 46532 40868 46560
rect 40543 46529 40555 46532
rect 40497 46523 40555 46529
rect 40862 46520 40868 46532
rect 40920 46520 40926 46572
rect 42242 46520 42248 46572
rect 42300 46560 42306 46572
rect 42720 46569 42748 46600
rect 42886 46588 42892 46600
rect 42944 46588 42950 46640
rect 43364 46628 43392 46656
rect 44726 46628 44732 46640
rect 43364 46600 43576 46628
rect 44687 46600 44732 46628
rect 42429 46563 42487 46569
rect 42429 46560 42441 46563
rect 42300 46532 42441 46560
rect 42300 46520 42306 46532
rect 42429 46529 42441 46532
rect 42475 46529 42487 46563
rect 42429 46523 42487 46529
rect 42705 46563 42763 46569
rect 42705 46529 42717 46563
rect 42751 46529 42763 46563
rect 42705 46523 42763 46529
rect 42794 46520 42800 46572
rect 42852 46560 42858 46572
rect 43548 46569 43576 46600
rect 44726 46588 44732 46600
rect 44784 46588 44790 46640
rect 44945 46631 45003 46637
rect 44945 46597 44957 46631
rect 44991 46628 45003 46631
rect 48682 46628 48688 46640
rect 44991 46600 48688 46628
rect 44991 46597 45003 46600
rect 44945 46591 45003 46597
rect 48682 46588 48688 46600
rect 48740 46588 48746 46640
rect 43349 46563 43407 46569
rect 43349 46560 43361 46563
rect 42852 46532 43361 46560
rect 42852 46520 42858 46532
rect 43349 46529 43361 46532
rect 43395 46529 43407 46563
rect 43349 46523 43407 46529
rect 43533 46563 43591 46569
rect 43533 46529 43545 46563
rect 43579 46529 43591 46563
rect 43533 46523 43591 46529
rect 43622 46520 43628 46572
rect 43680 46560 43686 46572
rect 43898 46560 43904 46572
rect 43680 46532 43725 46560
rect 43859 46532 43904 46560
rect 43680 46520 43686 46532
rect 43898 46520 43904 46532
rect 43956 46520 43962 46572
rect 45186 46520 45192 46572
rect 45244 46560 45250 46572
rect 45554 46560 45560 46572
rect 45244 46532 45560 46560
rect 45244 46520 45250 46532
rect 45554 46520 45560 46532
rect 45612 46520 45618 46572
rect 45738 46560 45744 46572
rect 45699 46532 45744 46560
rect 45738 46520 45744 46532
rect 45796 46520 45802 46572
rect 46842 46560 46848 46572
rect 46803 46532 46848 46560
rect 46842 46520 46848 46532
rect 46900 46520 46906 46572
rect 49786 46520 49792 46572
rect 49844 46560 49850 46572
rect 49881 46563 49939 46569
rect 49881 46560 49893 46563
rect 49844 46532 49893 46560
rect 49844 46520 49850 46532
rect 49881 46529 49893 46532
rect 49927 46529 49939 46563
rect 50062 46560 50068 46572
rect 50023 46532 50068 46560
rect 49881 46523 49939 46529
rect 50062 46520 50068 46532
rect 50120 46520 50126 46572
rect 50706 46560 50712 46572
rect 50667 46532 50712 46560
rect 50706 46520 50712 46532
rect 50764 46520 50770 46572
rect 56873 46563 56931 46569
rect 56873 46529 56885 46563
rect 56919 46529 56931 46563
rect 58066 46560 58072 46572
rect 58027 46532 58072 46560
rect 56873 46523 56931 46529
rect 40144 46492 40172 46520
rect 38120 46464 40172 46492
rect 41046 46452 41052 46504
rect 41104 46492 41110 46504
rect 43717 46495 43775 46501
rect 43717 46492 43729 46495
rect 41104 46464 43729 46492
rect 41104 46452 41110 46464
rect 43717 46461 43729 46464
rect 43763 46492 43775 46495
rect 44174 46492 44180 46504
rect 43763 46464 44180 46492
rect 43763 46461 43775 46464
rect 43717 46455 43775 46461
rect 44174 46452 44180 46464
rect 44232 46492 44238 46504
rect 45278 46492 45284 46504
rect 44232 46464 45284 46492
rect 44232 46452 44238 46464
rect 45278 46452 45284 46464
rect 45336 46452 45342 46504
rect 45649 46495 45707 46501
rect 45649 46461 45661 46495
rect 45695 46492 45707 46495
rect 46198 46492 46204 46504
rect 45695 46464 46204 46492
rect 45695 46461 45707 46464
rect 45649 46455 45707 46461
rect 46198 46452 46204 46464
rect 46256 46492 46262 46504
rect 46860 46492 46888 46520
rect 46256 46464 46888 46492
rect 47581 46495 47639 46501
rect 46256 46452 46262 46464
rect 47581 46461 47593 46495
rect 47627 46492 47639 46495
rect 47670 46492 47676 46504
rect 47627 46464 47676 46492
rect 47627 46461 47639 46464
rect 47581 46455 47639 46461
rect 47670 46452 47676 46464
rect 47728 46452 47734 46504
rect 47762 46452 47768 46504
rect 47820 46492 47826 46504
rect 47857 46495 47915 46501
rect 47857 46492 47869 46495
rect 47820 46464 47869 46492
rect 47820 46452 47826 46464
rect 47857 46461 47869 46464
rect 47903 46461 47915 46495
rect 47857 46455 47915 46461
rect 50801 46495 50859 46501
rect 50801 46461 50813 46495
rect 50847 46492 50859 46495
rect 51258 46492 51264 46504
rect 50847 46464 51264 46492
rect 50847 46461 50859 46464
rect 50801 46455 50859 46461
rect 51258 46452 51264 46464
rect 51316 46452 51322 46504
rect 38838 46384 38844 46436
rect 38896 46424 38902 46436
rect 39853 46427 39911 46433
rect 39853 46424 39865 46427
rect 38896 46396 39865 46424
rect 38896 46384 38902 46396
rect 39853 46393 39865 46396
rect 39899 46393 39911 46427
rect 56888 46424 56916 46523
rect 58066 46520 58072 46532
rect 58124 46520 58130 46572
rect 39853 46387 39911 46393
rect 41386 46396 56916 46424
rect 32442 46328 34468 46356
rect 36722 46316 36728 46368
rect 36780 46356 36786 46368
rect 38013 46359 38071 46365
rect 38013 46356 38025 46359
rect 36780 46328 38025 46356
rect 36780 46316 36786 46328
rect 38013 46325 38025 46328
rect 38059 46325 38071 46359
rect 38013 46319 38071 46325
rect 38470 46316 38476 46368
rect 38528 46356 38534 46368
rect 39209 46359 39267 46365
rect 39209 46356 39221 46359
rect 38528 46328 39221 46356
rect 38528 46316 38534 46328
rect 39209 46325 39221 46328
rect 39255 46325 39267 46359
rect 39209 46319 39267 46325
rect 39298 46316 39304 46368
rect 39356 46356 39362 46368
rect 41386 46356 41414 46396
rect 39356 46328 41414 46356
rect 42429 46359 42487 46365
rect 39356 46316 39362 46328
rect 42429 46325 42441 46359
rect 42475 46356 42487 46359
rect 42702 46356 42708 46368
rect 42475 46328 42708 46356
rect 42475 46325 42487 46328
rect 42429 46319 42487 46325
rect 42702 46316 42708 46328
rect 42760 46316 42766 46368
rect 44085 46359 44143 46365
rect 44085 46325 44097 46359
rect 44131 46356 44143 46359
rect 44913 46359 44971 46365
rect 44913 46356 44925 46359
rect 44131 46328 44925 46356
rect 44131 46325 44143 46328
rect 44085 46319 44143 46325
rect 44913 46325 44925 46328
rect 44959 46325 44971 46359
rect 44913 46319 44971 46325
rect 46937 46359 46995 46365
rect 46937 46325 46949 46359
rect 46983 46356 46995 46359
rect 48406 46356 48412 46368
rect 46983 46328 48412 46356
rect 46983 46325 46995 46328
rect 46937 46319 46995 46325
rect 48406 46316 48412 46328
rect 48464 46316 48470 46368
rect 49878 46356 49884 46368
rect 49791 46328 49884 46356
rect 49878 46316 49884 46328
rect 49936 46356 49942 46368
rect 50982 46356 50988 46368
rect 49936 46328 50988 46356
rect 49936 46316 49942 46328
rect 50982 46316 50988 46328
rect 51040 46316 51046 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 20530 46152 20536 46164
rect 18340 46124 20536 46152
rect 18340 46025 18368 46124
rect 20530 46112 20536 46124
rect 20588 46152 20594 46164
rect 20625 46155 20683 46161
rect 20625 46152 20637 46155
rect 20588 46124 20637 46152
rect 20588 46112 20594 46124
rect 20625 46121 20637 46124
rect 20671 46121 20683 46155
rect 20625 46115 20683 46121
rect 26050 46112 26056 46164
rect 26108 46152 26114 46164
rect 27065 46155 27123 46161
rect 27065 46152 27077 46155
rect 26108 46124 27077 46152
rect 26108 46112 26114 46124
rect 27065 46121 27077 46124
rect 27111 46152 27123 46155
rect 28994 46152 29000 46164
rect 27111 46124 28856 46152
rect 28955 46124 29000 46152
rect 27111 46121 27123 46124
rect 27065 46115 27123 46121
rect 20254 46044 20260 46096
rect 20312 46084 20318 46096
rect 21085 46087 21143 46093
rect 21085 46084 21097 46087
rect 20312 46056 21097 46084
rect 20312 46044 20318 46056
rect 21085 46053 21097 46056
rect 21131 46053 21143 46087
rect 21085 46047 21143 46053
rect 23109 46087 23167 46093
rect 23109 46053 23121 46087
rect 23155 46084 23167 46087
rect 23658 46084 23664 46096
rect 23155 46056 23664 46084
rect 23155 46053 23167 46056
rect 23109 46047 23167 46053
rect 23658 46044 23664 46056
rect 23716 46084 23722 46096
rect 24210 46084 24216 46096
rect 23716 46056 24216 46084
rect 23716 46044 23722 46056
rect 24210 46044 24216 46056
rect 24268 46044 24274 46096
rect 28828 46084 28856 46124
rect 28994 46112 29000 46124
rect 29052 46112 29058 46164
rect 33410 46152 33416 46164
rect 31036 46124 33416 46152
rect 31036 46084 31064 46124
rect 33410 46112 33416 46124
rect 33468 46152 33474 46164
rect 33468 46124 33640 46152
rect 33468 46112 33474 46124
rect 28828 46056 31064 46084
rect 33612 46084 33640 46124
rect 33686 46112 33692 46164
rect 33744 46152 33750 46164
rect 34793 46155 34851 46161
rect 34793 46152 34805 46155
rect 33744 46124 34805 46152
rect 33744 46112 33750 46124
rect 34793 46121 34805 46124
rect 34839 46121 34851 46155
rect 38378 46152 38384 46164
rect 34793 46115 34851 46121
rect 38028 46124 38384 46152
rect 35802 46084 35808 46096
rect 33612 46056 35808 46084
rect 18325 46019 18383 46025
rect 18325 45985 18337 46019
rect 18371 45985 18383 46019
rect 18325 45979 18383 45985
rect 18782 45976 18788 46028
rect 18840 46016 18846 46028
rect 19245 46019 19303 46025
rect 19245 46016 19257 46019
rect 18840 45988 19257 46016
rect 18840 45976 18846 45988
rect 19245 45985 19257 45988
rect 19291 45985 19303 46019
rect 21729 46019 21787 46025
rect 21729 46016 21741 46019
rect 19245 45979 19303 45985
rect 20272 45988 21741 46016
rect 18509 45951 18567 45957
rect 18509 45917 18521 45951
rect 18555 45948 18567 45951
rect 19150 45948 19156 45960
rect 18555 45920 19156 45948
rect 18555 45917 18567 45920
rect 18509 45911 18567 45917
rect 19150 45908 19156 45920
rect 19208 45908 19214 45960
rect 19260 45948 19288 45979
rect 20272 45948 20300 45988
rect 21729 45985 21741 45988
rect 21775 45985 21787 46019
rect 24394 46016 24400 46028
rect 21729 45979 21787 45985
rect 23492 45988 24400 46016
rect 21269 45951 21327 45957
rect 21269 45948 21281 45951
rect 19260 45920 20300 45948
rect 20364 45920 21281 45948
rect 19334 45840 19340 45892
rect 19392 45880 19398 45892
rect 19490 45883 19548 45889
rect 19490 45880 19502 45883
rect 19392 45852 19502 45880
rect 19392 45840 19398 45852
rect 19490 45849 19502 45852
rect 19536 45849 19548 45883
rect 19490 45843 19548 45849
rect 18693 45815 18751 45821
rect 18693 45781 18705 45815
rect 18739 45812 18751 45815
rect 20364 45812 20392 45920
rect 21269 45917 21281 45920
rect 21315 45917 21327 45951
rect 21744 45948 21772 45979
rect 22370 45948 22376 45960
rect 21744 45920 22376 45948
rect 21269 45911 21327 45917
rect 22370 45908 22376 45920
rect 22428 45948 22434 45960
rect 23106 45948 23112 45960
rect 22428 45920 23112 45948
rect 22428 45908 22434 45920
rect 23106 45908 23112 45920
rect 23164 45948 23170 45960
rect 23492 45948 23520 45988
rect 24394 45976 24400 45988
rect 24452 45976 24458 46028
rect 29730 45976 29736 46028
rect 29788 46016 29794 46028
rect 29917 46019 29975 46025
rect 29917 46016 29929 46019
rect 29788 45988 29929 46016
rect 29788 45976 29794 45988
rect 29917 45985 29929 45988
rect 29963 46016 29975 46019
rect 30374 46016 30380 46028
rect 29963 45988 30380 46016
rect 29963 45985 29975 45988
rect 29917 45979 29975 45985
rect 30374 45976 30380 45988
rect 30432 45976 30438 46028
rect 31018 46016 31024 46028
rect 30979 45988 31024 46016
rect 31018 45976 31024 45988
rect 31076 45976 31082 46028
rect 23164 45920 23520 45948
rect 23845 45951 23903 45957
rect 23164 45908 23170 45920
rect 23845 45917 23857 45951
rect 23891 45948 23903 45951
rect 24946 45948 24952 45960
rect 23891 45920 24952 45948
rect 23891 45917 23903 45920
rect 23845 45911 23903 45917
rect 24946 45908 24952 45920
rect 25004 45908 25010 45960
rect 27614 45948 27620 45960
rect 27575 45920 27620 45948
rect 27614 45908 27620 45920
rect 27672 45908 27678 45960
rect 28258 45908 28264 45960
rect 28316 45948 28322 45960
rect 29549 45951 29607 45957
rect 29549 45948 29561 45951
rect 28316 45920 29561 45948
rect 28316 45908 28322 45920
rect 29549 45917 29561 45920
rect 29595 45917 29607 45951
rect 29549 45911 29607 45917
rect 31288 45951 31346 45957
rect 31288 45917 31300 45951
rect 31334 45948 31346 45951
rect 32122 45948 32128 45960
rect 31334 45920 32128 45948
rect 31334 45917 31346 45920
rect 31288 45911 31346 45917
rect 32122 45908 32128 45920
rect 32180 45908 32186 45960
rect 33612 45957 33640 46056
rect 35802 46044 35808 46056
rect 35860 46044 35866 46096
rect 36265 46019 36323 46025
rect 36265 46016 36277 46019
rect 34900 45988 36277 46016
rect 34900 45960 34928 45988
rect 36265 45985 36277 45988
rect 36311 45985 36323 46019
rect 36265 45979 36323 45985
rect 33413 45951 33471 45957
rect 33413 45917 33425 45951
rect 33459 45917 33471 45951
rect 33413 45911 33471 45917
rect 33505 45951 33563 45957
rect 33505 45917 33517 45951
rect 33551 45917 33563 45951
rect 33505 45911 33563 45917
rect 33597 45951 33655 45957
rect 33597 45917 33609 45951
rect 33643 45917 33655 45951
rect 33778 45948 33784 45960
rect 33739 45920 33784 45948
rect 33597 45911 33655 45917
rect 21818 45840 21824 45892
rect 21876 45880 21882 45892
rect 24670 45889 24676 45892
rect 21974 45883 22032 45889
rect 21974 45880 21986 45883
rect 21876 45852 21986 45880
rect 21876 45840 21882 45852
rect 21974 45849 21986 45852
rect 22020 45849 22032 45883
rect 24664 45880 24676 45889
rect 21974 45843 22032 45849
rect 23676 45852 24676 45880
rect 23676 45821 23704 45852
rect 24664 45843 24676 45852
rect 24670 45840 24676 45843
rect 24728 45840 24734 45892
rect 26970 45880 26976 45892
rect 26931 45852 26976 45880
rect 26970 45840 26976 45852
rect 27028 45840 27034 45892
rect 27706 45840 27712 45892
rect 27764 45880 27770 45892
rect 27862 45883 27920 45889
rect 27862 45880 27874 45883
rect 27764 45852 27874 45880
rect 27764 45840 27770 45852
rect 27862 45849 27874 45852
rect 27908 45849 27920 45883
rect 27862 45843 27920 45849
rect 18739 45784 20392 45812
rect 23661 45815 23719 45821
rect 18739 45781 18751 45784
rect 18693 45775 18751 45781
rect 23661 45781 23673 45815
rect 23707 45781 23719 45815
rect 23661 45775 23719 45781
rect 25590 45772 25596 45824
rect 25648 45812 25654 45824
rect 25777 45815 25835 45821
rect 25777 45812 25789 45815
rect 25648 45784 25789 45812
rect 25648 45772 25654 45784
rect 25777 45781 25789 45784
rect 25823 45781 25835 45815
rect 25777 45775 25835 45781
rect 32401 45815 32459 45821
rect 32401 45781 32413 45815
rect 32447 45812 32459 45815
rect 32582 45812 32588 45824
rect 32447 45784 32588 45812
rect 32447 45781 32459 45784
rect 32401 45775 32459 45781
rect 32582 45772 32588 45784
rect 32640 45772 32646 45824
rect 33134 45812 33140 45824
rect 33095 45784 33140 45812
rect 33134 45772 33140 45784
rect 33192 45772 33198 45824
rect 33428 45812 33456 45911
rect 33520 45880 33548 45911
rect 33778 45908 33784 45920
rect 33836 45908 33842 45960
rect 34701 45951 34759 45957
rect 34701 45917 34713 45951
rect 34747 45917 34759 45951
rect 34882 45948 34888 45960
rect 34843 45920 34888 45948
rect 34701 45911 34759 45917
rect 33686 45880 33692 45892
rect 33520 45852 33692 45880
rect 33686 45840 33692 45852
rect 33744 45840 33750 45892
rect 34716 45880 34744 45911
rect 34882 45908 34888 45920
rect 34940 45908 34946 45960
rect 35986 45948 35992 45960
rect 35947 45920 35992 45948
rect 35986 45908 35992 45920
rect 36044 45908 36050 45960
rect 36081 45951 36139 45957
rect 36081 45917 36093 45951
rect 36127 45948 36139 45951
rect 36998 45948 37004 45960
rect 36127 45920 37004 45948
rect 36127 45917 36139 45920
rect 36081 45911 36139 45917
rect 36998 45908 37004 45920
rect 37056 45908 37062 45960
rect 37645 45951 37703 45957
rect 37645 45917 37657 45951
rect 37691 45948 37703 45951
rect 37826 45948 37832 45960
rect 37691 45920 37832 45948
rect 37691 45917 37703 45920
rect 37645 45911 37703 45917
rect 37826 45908 37832 45920
rect 37884 45908 37890 45960
rect 37921 45951 37979 45957
rect 37921 45917 37933 45951
rect 37967 45948 37979 45951
rect 38028 45948 38056 46124
rect 38378 46112 38384 46124
rect 38436 46152 38442 46164
rect 42702 46152 42708 46164
rect 38436 46124 42708 46152
rect 38436 46112 38442 46124
rect 42702 46112 42708 46124
rect 42760 46112 42766 46164
rect 45002 46112 45008 46164
rect 45060 46152 45066 46164
rect 45097 46155 45155 46161
rect 45097 46152 45109 46155
rect 45060 46124 45109 46152
rect 45060 46112 45066 46124
rect 45097 46121 45109 46124
rect 45143 46121 45155 46155
rect 45097 46115 45155 46121
rect 45649 46155 45707 46161
rect 45649 46121 45661 46155
rect 45695 46152 45707 46155
rect 45738 46152 45744 46164
rect 45695 46124 45744 46152
rect 45695 46121 45707 46124
rect 45649 46115 45707 46121
rect 45738 46112 45744 46124
rect 45796 46112 45802 46164
rect 47762 46152 47768 46164
rect 47723 46124 47768 46152
rect 47762 46112 47768 46124
rect 47820 46112 47826 46164
rect 47946 46152 47952 46164
rect 47907 46124 47952 46152
rect 47946 46112 47952 46124
rect 48004 46112 48010 46164
rect 38580 46056 40356 46084
rect 37967 45920 38056 45948
rect 37967 45917 37979 45920
rect 37921 45911 37979 45917
rect 38102 45908 38108 45960
rect 38160 45948 38166 45960
rect 38160 45920 38205 45948
rect 38160 45908 38166 45920
rect 38470 45908 38476 45960
rect 38528 45948 38534 45960
rect 38580 45957 38608 46056
rect 39114 45976 39120 46028
rect 39172 46016 39178 46028
rect 39172 45988 40264 46016
rect 39172 45976 39178 45988
rect 38565 45951 38623 45957
rect 38565 45948 38577 45951
rect 38528 45920 38577 45948
rect 38528 45908 38534 45920
rect 38565 45917 38577 45920
rect 38611 45917 38623 45951
rect 38930 45948 38936 45960
rect 38891 45920 38936 45948
rect 38565 45911 38623 45917
rect 38930 45908 38936 45920
rect 38988 45908 38994 45960
rect 40236 45957 40264 45988
rect 40328 45957 40356 46056
rect 41230 46044 41236 46096
rect 41288 46084 41294 46096
rect 43162 46084 43168 46096
rect 41288 46056 43168 46084
rect 41288 46044 41294 46056
rect 43162 46044 43168 46056
rect 43220 46044 43226 46096
rect 45554 46044 45560 46096
rect 45612 46084 45618 46096
rect 49878 46084 49884 46096
rect 45612 46056 49884 46084
rect 45612 46044 45618 46056
rect 49878 46044 49884 46056
rect 49936 46044 49942 46096
rect 42886 46016 42892 46028
rect 42352 45988 42892 46016
rect 40129 45951 40187 45957
rect 40129 45917 40141 45951
rect 40175 45917 40187 45951
rect 40129 45911 40187 45917
rect 40221 45951 40279 45957
rect 40221 45917 40233 45951
rect 40267 45917 40279 45951
rect 40221 45911 40279 45917
rect 40313 45951 40371 45957
rect 40313 45917 40325 45951
rect 40359 45917 40371 45951
rect 40313 45911 40371 45917
rect 40497 45951 40555 45957
rect 40497 45917 40509 45951
rect 40543 45948 40555 45951
rect 41049 45951 41107 45957
rect 41049 45948 41061 45951
rect 40543 45920 41061 45948
rect 40543 45917 40555 45920
rect 40497 45911 40555 45917
rect 41049 45917 41061 45920
rect 41095 45917 41107 45951
rect 41049 45911 41107 45917
rect 41233 45951 41291 45957
rect 41233 45917 41245 45951
rect 41279 45948 41291 45951
rect 41690 45948 41696 45960
rect 41279 45920 41696 45948
rect 41279 45917 41291 45920
rect 41233 45911 41291 45917
rect 37182 45880 37188 45892
rect 34716 45852 37188 45880
rect 37182 45840 37188 45852
rect 37240 45840 37246 45892
rect 38746 45880 38752 45892
rect 38707 45852 38752 45880
rect 38746 45840 38752 45852
rect 38804 45840 38810 45892
rect 38841 45883 38899 45889
rect 38841 45849 38853 45883
rect 38887 45880 38899 45883
rect 40034 45880 40040 45892
rect 38887 45852 40040 45880
rect 38887 45849 38899 45852
rect 38841 45843 38899 45849
rect 40034 45840 40040 45852
rect 40092 45840 40098 45892
rect 40144 45880 40172 45911
rect 40770 45880 40776 45892
rect 40144 45852 40776 45880
rect 40770 45840 40776 45852
rect 40828 45840 40834 45892
rect 41064 45880 41092 45911
rect 41690 45908 41696 45920
rect 41748 45908 41754 45960
rect 42352 45957 42380 45988
rect 42886 45976 42892 45988
rect 42944 45976 42950 46028
rect 43898 45976 43904 46028
rect 43956 46016 43962 46028
rect 43956 45988 45876 46016
rect 43956 45976 43962 45988
rect 42337 45951 42395 45957
rect 42337 45917 42349 45951
rect 42383 45917 42395 45951
rect 42702 45948 42708 45960
rect 42663 45920 42708 45948
rect 42337 45911 42395 45917
rect 42702 45908 42708 45920
rect 42760 45908 42766 45960
rect 42794 45908 42800 45960
rect 42852 45948 42858 45960
rect 42852 45920 42897 45948
rect 42852 45908 42858 45920
rect 42978 45908 42984 45960
rect 43036 45948 43042 45960
rect 43622 45948 43628 45960
rect 43036 45920 43628 45948
rect 43036 45908 43042 45920
rect 43622 45908 43628 45920
rect 43680 45908 43686 45960
rect 44174 45948 44180 45960
rect 44135 45920 44180 45948
rect 44174 45908 44180 45920
rect 44232 45908 44238 45960
rect 44450 45908 44456 45960
rect 44508 45948 44514 45960
rect 44910 45948 44916 45960
rect 44508 45920 44916 45948
rect 44508 45908 44514 45920
rect 44910 45908 44916 45920
rect 44968 45948 44974 45960
rect 45848 45957 45876 45988
rect 45005 45951 45063 45957
rect 45005 45948 45017 45951
rect 44968 45920 45017 45948
rect 44968 45908 44974 45920
rect 45005 45917 45017 45920
rect 45051 45917 45063 45951
rect 45005 45911 45063 45917
rect 45189 45951 45247 45957
rect 45189 45917 45201 45951
rect 45235 45917 45247 45951
rect 45189 45911 45247 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45917 45707 45951
rect 45649 45911 45707 45917
rect 45833 45951 45891 45957
rect 45833 45917 45845 45951
rect 45879 45948 45891 45951
rect 50154 45948 50160 45960
rect 45879 45920 50160 45948
rect 45879 45917 45891 45920
rect 45833 45911 45891 45917
rect 41064 45852 41414 45880
rect 35526 45812 35532 45824
rect 33428 45784 35532 45812
rect 35526 45772 35532 45784
rect 35584 45772 35590 45824
rect 36262 45812 36268 45824
rect 36223 45784 36268 45812
rect 36262 45772 36268 45784
rect 36320 45772 36326 45824
rect 36630 45772 36636 45824
rect 36688 45812 36694 45824
rect 37734 45812 37740 45824
rect 36688 45784 37740 45812
rect 36688 45772 36694 45784
rect 37734 45772 37740 45784
rect 37792 45812 37798 45824
rect 37829 45815 37887 45821
rect 37829 45812 37841 45815
rect 37792 45784 37841 45812
rect 37792 45772 37798 45784
rect 37829 45781 37841 45784
rect 37875 45781 37887 45815
rect 37829 45775 37887 45781
rect 37918 45772 37924 45824
rect 37976 45812 37982 45824
rect 39117 45815 39175 45821
rect 39117 45812 39129 45815
rect 37976 45784 39129 45812
rect 37976 45772 37982 45784
rect 39117 45781 39129 45784
rect 39163 45781 39175 45815
rect 39850 45812 39856 45824
rect 39811 45784 39856 45812
rect 39117 45775 39175 45781
rect 39850 45772 39856 45784
rect 39908 45772 39914 45824
rect 40494 45772 40500 45824
rect 40552 45812 40558 45824
rect 41141 45815 41199 45821
rect 41141 45812 41153 45815
rect 40552 45784 41153 45812
rect 40552 45772 40558 45784
rect 41141 45781 41153 45784
rect 41187 45781 41199 45815
rect 41386 45812 41414 45852
rect 42242 45840 42248 45892
rect 42300 45880 42306 45892
rect 42429 45883 42487 45889
rect 42429 45880 42441 45883
rect 42300 45852 42441 45880
rect 42300 45840 42306 45852
rect 42429 45849 42441 45852
rect 42475 45849 42487 45883
rect 42429 45843 42487 45849
rect 42521 45883 42579 45889
rect 42521 45849 42533 45883
rect 42567 45880 42579 45883
rect 43346 45880 43352 45892
rect 42567 45852 43352 45880
rect 42567 45849 42579 45852
rect 42521 45843 42579 45849
rect 43346 45840 43352 45852
rect 43404 45840 43410 45892
rect 44542 45840 44548 45892
rect 44600 45880 44606 45892
rect 45204 45880 45232 45911
rect 44600 45852 45232 45880
rect 45664 45880 45692 45911
rect 50154 45908 50160 45920
rect 50212 45908 50218 45960
rect 50982 45948 50988 45960
rect 50943 45920 50988 45948
rect 50982 45908 50988 45920
rect 51040 45908 51046 45960
rect 51258 45948 51264 45960
rect 51171 45920 51264 45948
rect 51258 45908 51264 45920
rect 51316 45948 51322 45960
rect 51810 45948 51816 45960
rect 51316 45920 51816 45948
rect 51316 45908 51322 45920
rect 51810 45908 51816 45920
rect 51868 45908 51874 45960
rect 56870 45908 56876 45960
rect 56928 45948 56934 45960
rect 56965 45951 57023 45957
rect 56965 45948 56977 45951
rect 56928 45920 56977 45948
rect 56928 45908 56934 45920
rect 56965 45917 56977 45920
rect 57011 45948 57023 45951
rect 57422 45948 57428 45960
rect 57011 45920 57428 45948
rect 57011 45917 57023 45920
rect 56965 45911 57023 45917
rect 57422 45908 57428 45920
rect 57480 45908 57486 45960
rect 57790 45948 57796 45960
rect 57751 45920 57796 45948
rect 57790 45908 57796 45920
rect 57848 45908 57854 45960
rect 46290 45880 46296 45892
rect 45664 45852 46296 45880
rect 44600 45840 44606 45852
rect 46290 45840 46296 45852
rect 46348 45840 46354 45892
rect 47118 45840 47124 45892
rect 47176 45880 47182 45892
rect 47578 45880 47584 45892
rect 47176 45852 47584 45880
rect 47176 45840 47182 45852
rect 47578 45840 47584 45852
rect 47636 45840 47642 45892
rect 50801 45883 50859 45889
rect 50801 45849 50813 45883
rect 50847 45880 50859 45883
rect 52086 45880 52092 45892
rect 50847 45852 52092 45880
rect 50847 45849 50859 45852
rect 50801 45843 50859 45849
rect 52086 45840 52092 45852
rect 52144 45840 52150 45892
rect 41690 45812 41696 45824
rect 41386 45784 41696 45812
rect 41141 45775 41199 45781
rect 41690 45772 41696 45784
rect 41748 45772 41754 45824
rect 42150 45812 42156 45824
rect 42111 45784 42156 45812
rect 42150 45772 42156 45784
rect 42208 45772 42214 45824
rect 43070 45772 43076 45824
rect 43128 45812 43134 45824
rect 44269 45815 44327 45821
rect 44269 45812 44281 45815
rect 43128 45784 44281 45812
rect 43128 45772 43134 45784
rect 44269 45781 44281 45784
rect 44315 45781 44327 45815
rect 44269 45775 44327 45781
rect 45002 45772 45008 45824
rect 45060 45812 45066 45824
rect 45646 45812 45652 45824
rect 45060 45784 45652 45812
rect 45060 45772 45066 45784
rect 45646 45772 45652 45784
rect 45704 45772 45710 45824
rect 47210 45772 47216 45824
rect 47268 45812 47274 45824
rect 47781 45815 47839 45821
rect 47781 45812 47793 45815
rect 47268 45784 47793 45812
rect 47268 45772 47274 45784
rect 47781 45781 47793 45784
rect 47827 45812 47839 45815
rect 47946 45812 47952 45824
rect 47827 45784 47952 45812
rect 47827 45781 47839 45784
rect 47781 45775 47839 45781
rect 47946 45772 47952 45784
rect 48004 45772 48010 45824
rect 50706 45772 50712 45824
rect 50764 45812 50770 45824
rect 51169 45815 51227 45821
rect 51169 45812 51181 45815
rect 50764 45784 51181 45812
rect 50764 45772 50770 45784
rect 51169 45781 51181 45784
rect 51215 45781 51227 45815
rect 57054 45812 57060 45824
rect 57015 45784 57060 45812
rect 51169 45775 51227 45781
rect 57054 45772 57060 45784
rect 57112 45772 57118 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 20438 45568 20444 45620
rect 20496 45608 20502 45620
rect 20993 45611 21051 45617
rect 20993 45608 21005 45611
rect 20496 45580 21005 45608
rect 20496 45568 20502 45580
rect 20993 45577 21005 45580
rect 21039 45577 21051 45611
rect 20993 45571 21051 45577
rect 24964 45580 26372 45608
rect 2038 45500 2044 45552
rect 2096 45540 2102 45552
rect 22646 45549 22652 45552
rect 22640 45540 22652 45549
rect 2096 45512 22508 45540
rect 22607 45512 22652 45540
rect 2096 45500 2102 45512
rect 18782 45432 18788 45484
rect 18840 45472 18846 45484
rect 18877 45475 18935 45481
rect 18877 45472 18889 45475
rect 18840 45444 18889 45472
rect 18840 45432 18846 45444
rect 18877 45441 18889 45444
rect 18923 45441 18935 45475
rect 18877 45435 18935 45441
rect 19144 45475 19202 45481
rect 19144 45441 19156 45475
rect 19190 45472 19202 45475
rect 20254 45472 20260 45484
rect 19190 45444 20260 45472
rect 19190 45441 19202 45444
rect 19144 45435 19202 45441
rect 20254 45432 20260 45444
rect 20312 45432 20318 45484
rect 20530 45432 20536 45484
rect 20588 45472 20594 45484
rect 20717 45475 20775 45481
rect 20717 45472 20729 45475
rect 20588 45444 20729 45472
rect 20588 45432 20594 45444
rect 20717 45441 20729 45444
rect 20763 45441 20775 45475
rect 20717 45435 20775 45441
rect 20901 45475 20959 45481
rect 20901 45441 20913 45475
rect 20947 45441 20959 45475
rect 20901 45435 20959 45441
rect 21085 45475 21143 45481
rect 21085 45441 21097 45475
rect 21131 45441 21143 45475
rect 21085 45435 21143 45441
rect 21269 45475 21327 45481
rect 21269 45441 21281 45475
rect 21315 45472 21327 45475
rect 22094 45472 22100 45484
rect 21315 45444 22100 45472
rect 21315 45441 21327 45444
rect 21269 45435 21327 45441
rect 20162 45296 20168 45348
rect 20220 45336 20226 45348
rect 20916 45336 20944 45435
rect 20220 45308 20944 45336
rect 20220 45296 20226 45308
rect 20257 45271 20315 45277
rect 20257 45237 20269 45271
rect 20303 45268 20315 45271
rect 20346 45268 20352 45280
rect 20303 45240 20352 45268
rect 20303 45237 20315 45240
rect 20257 45231 20315 45237
rect 20346 45228 20352 45240
rect 20404 45268 20410 45280
rect 21100 45268 21128 45435
rect 22094 45432 22100 45444
rect 22152 45432 22158 45484
rect 22480 45472 22508 45512
rect 22640 45503 22652 45512
rect 22646 45500 22652 45503
rect 22704 45500 22710 45552
rect 24964 45540 24992 45580
rect 25130 45540 25136 45552
rect 23676 45512 24992 45540
rect 25091 45512 25136 45540
rect 23676 45472 23704 45512
rect 25130 45500 25136 45512
rect 25188 45500 25194 45552
rect 25590 45500 25596 45552
rect 25648 45540 25654 45552
rect 26344 45540 26372 45580
rect 33778 45568 33784 45620
rect 33836 45608 33842 45620
rect 34425 45611 34483 45617
rect 34425 45608 34437 45611
rect 33836 45580 34437 45608
rect 33836 45568 33842 45580
rect 34425 45577 34437 45580
rect 34471 45577 34483 45611
rect 37918 45608 37924 45620
rect 34425 45571 34483 45577
rect 34992 45580 37924 45608
rect 27341 45543 27399 45549
rect 27341 45540 27353 45543
rect 25648 45512 26280 45540
rect 26344 45512 27353 45540
rect 25648 45500 25654 45512
rect 25682 45472 25688 45484
rect 22480 45444 23704 45472
rect 23768 45444 25688 45472
rect 22370 45404 22376 45416
rect 22331 45376 22376 45404
rect 22370 45364 22376 45376
rect 22428 45364 22434 45416
rect 23768 45345 23796 45444
rect 25682 45432 25688 45444
rect 25740 45472 25746 45484
rect 26252 45481 26280 45512
rect 27341 45509 27353 45512
rect 27387 45540 27399 45543
rect 27985 45543 28043 45549
rect 27985 45540 27997 45543
rect 27387 45512 27997 45540
rect 27387 45509 27399 45512
rect 27341 45503 27399 45509
rect 27985 45509 27997 45512
rect 28031 45540 28043 45543
rect 28442 45540 28448 45552
rect 28031 45512 28448 45540
rect 28031 45509 28043 45512
rect 27985 45503 28043 45509
rect 28442 45500 28448 45512
rect 28500 45500 28506 45552
rect 30006 45500 30012 45552
rect 30064 45540 30070 45552
rect 30101 45543 30159 45549
rect 30101 45540 30113 45543
rect 30064 45512 30113 45540
rect 30064 45500 30070 45512
rect 30101 45509 30113 45512
rect 30147 45509 30159 45543
rect 30101 45503 30159 45509
rect 32392 45543 32450 45549
rect 32392 45509 32404 45543
rect 32438 45540 32450 45543
rect 33134 45540 33140 45552
rect 32438 45512 33140 45540
rect 32438 45509 32450 45512
rect 32392 45503 32450 45509
rect 33134 45500 33140 45512
rect 33192 45500 33198 45552
rect 34992 45540 35020 45580
rect 37918 45568 37924 45580
rect 37976 45568 37982 45620
rect 38746 45568 38752 45620
rect 38804 45608 38810 45620
rect 38933 45611 38991 45617
rect 38933 45608 38945 45611
rect 38804 45580 38945 45608
rect 38804 45568 38810 45580
rect 38933 45577 38945 45580
rect 38979 45577 38991 45611
rect 38933 45571 38991 45577
rect 39850 45568 39856 45620
rect 39908 45608 39914 45620
rect 39908 45580 41828 45608
rect 39908 45568 39914 45580
rect 39942 45540 39948 45552
rect 34348 45512 35020 45540
rect 35268 45512 39948 45540
rect 26053 45475 26111 45481
rect 26053 45472 26065 45475
rect 25740 45444 26065 45472
rect 25740 45432 25746 45444
rect 26053 45441 26065 45444
rect 26099 45441 26111 45475
rect 26053 45435 26111 45441
rect 26237 45475 26295 45481
rect 26237 45441 26249 45475
rect 26283 45441 26295 45475
rect 26237 45435 26295 45441
rect 27709 45475 27767 45481
rect 27709 45441 27721 45475
rect 27755 45472 27767 45475
rect 28258 45472 28264 45484
rect 27755 45444 28264 45472
rect 27755 45441 27767 45444
rect 27709 45435 27767 45441
rect 28258 45432 28264 45444
rect 28316 45432 28322 45484
rect 34348 45481 34376 45512
rect 34333 45475 34391 45481
rect 34333 45441 34345 45475
rect 34379 45441 34391 45475
rect 34333 45435 34391 45441
rect 34517 45475 34575 45481
rect 34517 45441 34529 45475
rect 34563 45472 34575 45475
rect 34882 45472 34888 45484
rect 34563 45444 34888 45472
rect 34563 45441 34575 45444
rect 34517 45435 34575 45441
rect 34882 45432 34888 45444
rect 34940 45432 34946 45484
rect 34977 45475 35035 45481
rect 34977 45441 34989 45475
rect 35023 45441 35035 45475
rect 34977 45435 35035 45441
rect 35161 45475 35219 45481
rect 35161 45441 35173 45475
rect 35207 45474 35219 45475
rect 35268 45474 35296 45512
rect 39942 45500 39948 45512
rect 40000 45500 40006 45552
rect 40034 45500 40040 45552
rect 40092 45540 40098 45552
rect 40221 45543 40279 45549
rect 40221 45540 40233 45543
rect 40092 45512 40233 45540
rect 40092 45500 40098 45512
rect 40221 45509 40233 45512
rect 40267 45509 40279 45543
rect 40221 45503 40279 45509
rect 35207 45446 35296 45474
rect 35345 45475 35403 45481
rect 35207 45441 35219 45446
rect 35161 45435 35219 45441
rect 35345 45441 35357 45475
rect 35391 45441 35403 45475
rect 35345 45435 35403 45441
rect 35529 45475 35587 45481
rect 35529 45441 35541 45475
rect 35575 45472 35587 45475
rect 35618 45472 35624 45484
rect 35575 45444 35624 45472
rect 35575 45441 35587 45444
rect 35529 45435 35587 45441
rect 24210 45404 24216 45416
rect 24123 45376 24216 45404
rect 24210 45364 24216 45376
rect 24268 45404 24274 45416
rect 28994 45404 29000 45416
rect 24268 45376 25452 45404
rect 28955 45376 29000 45404
rect 24268 45364 24274 45376
rect 23753 45339 23811 45345
rect 23753 45305 23765 45339
rect 23799 45305 23811 45339
rect 23753 45299 23811 45305
rect 24581 45339 24639 45345
rect 24581 45305 24593 45339
rect 24627 45336 24639 45339
rect 25130 45336 25136 45348
rect 24627 45308 25136 45336
rect 24627 45305 24639 45308
rect 24581 45299 24639 45305
rect 25130 45296 25136 45308
rect 25188 45296 25194 45348
rect 25424 45345 25452 45376
rect 28994 45364 29000 45376
rect 29052 45364 29058 45416
rect 31018 45364 31024 45416
rect 31076 45404 31082 45416
rect 32125 45407 32183 45413
rect 32125 45404 32137 45407
rect 31076 45376 32137 45404
rect 31076 45364 31082 45376
rect 32125 45373 32137 45376
rect 32171 45373 32183 45407
rect 32125 45367 32183 45373
rect 25409 45339 25467 45345
rect 25409 45305 25421 45339
rect 25455 45305 25467 45339
rect 25409 45299 25467 45305
rect 30285 45339 30343 45345
rect 30285 45305 30297 45339
rect 30331 45336 30343 45339
rect 32030 45336 32036 45348
rect 30331 45308 32036 45336
rect 30331 45305 30343 45308
rect 30285 45299 30343 45305
rect 32030 45296 32036 45308
rect 32088 45296 32094 45348
rect 24670 45268 24676 45280
rect 20404 45240 21128 45268
rect 24631 45240 24676 45268
rect 20404 45228 20410 45240
rect 24670 45228 24676 45240
rect 24728 45228 24734 45280
rect 24762 45228 24768 45280
rect 24820 45268 24826 45280
rect 25593 45271 25651 45277
rect 25593 45268 25605 45271
rect 24820 45240 25605 45268
rect 24820 45228 24826 45240
rect 25593 45237 25605 45240
rect 25639 45237 25651 45271
rect 26050 45268 26056 45280
rect 26011 45240 26056 45268
rect 25593 45231 25651 45237
rect 26050 45228 26056 45240
rect 26108 45228 26114 45280
rect 32140 45268 32168 45367
rect 34606 45364 34612 45416
rect 34664 45404 34670 45416
rect 34992 45404 35020 45435
rect 35253 45407 35311 45413
rect 35253 45404 35265 45407
rect 34664 45376 35020 45404
rect 35176 45376 35265 45404
rect 34664 45364 34670 45376
rect 33410 45268 33416 45280
rect 32140 45240 33416 45268
rect 33410 45228 33416 45240
rect 33468 45228 33474 45280
rect 33505 45271 33563 45277
rect 33505 45237 33517 45271
rect 33551 45268 33563 45271
rect 33686 45268 33692 45280
rect 33551 45240 33692 45268
rect 33551 45237 33563 45240
rect 33505 45231 33563 45237
rect 33686 45228 33692 45240
rect 33744 45228 33750 45280
rect 35176 45268 35204 45376
rect 35253 45373 35265 45376
rect 35299 45373 35311 45407
rect 35360 45404 35388 45435
rect 35618 45432 35624 45444
rect 35676 45432 35682 45484
rect 36446 45472 36452 45484
rect 36407 45444 36452 45472
rect 36446 45432 36452 45444
rect 36504 45432 36510 45484
rect 36630 45472 36636 45484
rect 36591 45444 36636 45472
rect 36630 45432 36636 45444
rect 36688 45432 36694 45484
rect 36722 45432 36728 45484
rect 36780 45472 36786 45484
rect 37553 45475 37611 45481
rect 37553 45474 37565 45475
rect 37476 45472 37565 45474
rect 36780 45446 37565 45472
rect 36780 45444 37504 45446
rect 36780 45432 36786 45444
rect 37553 45441 37565 45446
rect 37599 45441 37611 45475
rect 37734 45472 37740 45484
rect 37695 45444 37740 45472
rect 37553 45435 37611 45441
rect 37734 45432 37740 45444
rect 37792 45432 37798 45484
rect 37830 45475 37888 45481
rect 37830 45441 37842 45475
rect 37876 45474 37888 45475
rect 37876 45472 38056 45474
rect 38286 45472 38292 45484
rect 37876 45446 38292 45472
rect 37876 45441 37888 45446
rect 38028 45444 38292 45446
rect 37830 45435 37888 45441
rect 38286 45432 38292 45444
rect 38344 45432 38350 45484
rect 38562 45472 38568 45484
rect 38523 45444 38568 45472
rect 38562 45432 38568 45444
rect 38620 45432 38626 45484
rect 39758 45432 39764 45484
rect 39816 45472 39822 45484
rect 40405 45475 40463 45481
rect 40405 45472 40417 45475
rect 39816 45444 40417 45472
rect 39816 45432 39822 45444
rect 40405 45441 40417 45444
rect 40451 45441 40463 45475
rect 40405 45435 40463 45441
rect 40494 45432 40500 45484
rect 40552 45472 40558 45484
rect 40681 45475 40739 45481
rect 40552 45444 40597 45472
rect 40552 45432 40558 45444
rect 40681 45441 40693 45475
rect 40727 45441 40739 45475
rect 40681 45435 40739 45441
rect 40865 45475 40923 45481
rect 40865 45441 40877 45475
rect 40911 45441 40923 45475
rect 40865 45435 40923 45441
rect 37634 45407 37692 45413
rect 35360 45376 35664 45404
rect 35253 45367 35311 45373
rect 35636 45348 35664 45376
rect 37634 45373 37646 45407
rect 37680 45404 37692 45407
rect 38657 45407 38715 45413
rect 37680 45376 37872 45404
rect 37680 45373 37692 45376
rect 37634 45367 37692 45373
rect 35618 45296 35624 45348
rect 35676 45296 35682 45348
rect 37844 45336 37872 45376
rect 38657 45373 38669 45407
rect 38703 45404 38715 45407
rect 39114 45404 39120 45416
rect 38703 45376 39120 45404
rect 38703 45373 38715 45376
rect 38657 45367 38715 45373
rect 39114 45364 39120 45376
rect 39172 45364 39178 45416
rect 40696 45404 40724 45435
rect 40512 45376 40724 45404
rect 40512 45348 40540 45376
rect 37918 45336 37924 45348
rect 37844 45308 37924 45336
rect 37918 45296 37924 45308
rect 37976 45296 37982 45348
rect 38010 45296 38016 45348
rect 38068 45336 38074 45348
rect 38068 45308 38792 45336
rect 38068 45296 38074 45308
rect 35434 45268 35440 45280
rect 35176 45240 35440 45268
rect 35434 45228 35440 45240
rect 35492 45228 35498 45280
rect 35710 45268 35716 45280
rect 35671 45240 35716 45268
rect 35710 45228 35716 45240
rect 35768 45228 35774 45280
rect 35986 45228 35992 45280
rect 36044 45268 36050 45280
rect 36446 45268 36452 45280
rect 36044 45240 36452 45268
rect 36044 45228 36050 45240
rect 36446 45228 36452 45240
rect 36504 45228 36510 45280
rect 36998 45228 37004 45280
rect 37056 45268 37062 45280
rect 37369 45271 37427 45277
rect 37369 45268 37381 45271
rect 37056 45240 37381 45268
rect 37056 45228 37062 45240
rect 37369 45237 37381 45240
rect 37415 45237 37427 45271
rect 37369 45231 37427 45237
rect 38194 45228 38200 45280
rect 38252 45268 38258 45280
rect 38654 45268 38660 45280
rect 38252 45240 38660 45268
rect 38252 45228 38258 45240
rect 38654 45228 38660 45240
rect 38712 45228 38718 45280
rect 38764 45268 38792 45308
rect 40494 45296 40500 45348
rect 40552 45296 40558 45348
rect 40589 45339 40647 45345
rect 40589 45305 40601 45339
rect 40635 45336 40647 45339
rect 40770 45336 40776 45348
rect 40635 45308 40776 45336
rect 40635 45305 40647 45308
rect 40589 45299 40647 45305
rect 40770 45296 40776 45308
rect 40828 45296 40834 45348
rect 40880 45336 40908 45435
rect 41230 45432 41236 45484
rect 41288 45472 41294 45484
rect 41800 45481 41828 45580
rect 42058 45568 42064 45620
rect 42116 45608 42122 45620
rect 42116 45580 43035 45608
rect 42116 45568 42122 45580
rect 42794 45540 42800 45552
rect 42444 45512 42800 45540
rect 42444 45481 42472 45512
rect 42794 45500 42800 45512
rect 42852 45500 42858 45552
rect 41693 45475 41751 45481
rect 41693 45472 41705 45475
rect 41288 45444 41705 45472
rect 41288 45432 41294 45444
rect 41693 45441 41705 45444
rect 41739 45441 41751 45475
rect 41693 45435 41751 45441
rect 41785 45475 41843 45481
rect 41785 45441 41797 45475
rect 41831 45441 41843 45475
rect 41785 45435 41843 45441
rect 42429 45475 42487 45481
rect 42429 45441 42441 45475
rect 42475 45441 42487 45475
rect 42429 45435 42487 45441
rect 42613 45475 42671 45481
rect 42613 45441 42625 45475
rect 42659 45441 42671 45475
rect 42613 45435 42671 45441
rect 42705 45475 42763 45481
rect 42705 45441 42717 45475
rect 42751 45472 42763 45475
rect 42886 45472 42892 45484
rect 42751 45444 42892 45472
rect 42751 45441 42763 45444
rect 42705 45435 42763 45441
rect 40954 45364 40960 45416
rect 41012 45404 41018 45416
rect 41509 45407 41567 45413
rect 41509 45404 41521 45407
rect 41012 45376 41521 45404
rect 41012 45364 41018 45376
rect 41509 45373 41521 45376
rect 41555 45373 41567 45407
rect 41509 45367 41567 45373
rect 41598 45364 41604 45416
rect 41656 45404 41662 45416
rect 41656 45376 41701 45404
rect 41656 45364 41662 45376
rect 41874 45364 41880 45416
rect 41932 45404 41938 45416
rect 42628 45404 42656 45435
rect 42886 45432 42892 45444
rect 42944 45432 42950 45484
rect 43007 45481 43035 45580
rect 43438 45568 43444 45620
rect 43496 45608 43502 45620
rect 48041 45611 48099 45617
rect 48041 45608 48053 45611
rect 43496 45580 48053 45608
rect 43496 45568 43502 45580
rect 48041 45577 48053 45580
rect 48087 45577 48099 45611
rect 48041 45571 48099 45577
rect 43162 45500 43168 45552
rect 43220 45540 43226 45552
rect 45741 45543 45799 45549
rect 45741 45540 45753 45543
rect 43220 45512 45753 45540
rect 43220 45500 43226 45512
rect 45741 45509 45753 45512
rect 45787 45540 45799 45543
rect 45830 45540 45836 45552
rect 45787 45512 45836 45540
rect 45787 45509 45799 45512
rect 45741 45503 45799 45509
rect 45830 45500 45836 45512
rect 45888 45500 45894 45552
rect 48774 45500 48780 45552
rect 48832 45540 48838 45552
rect 49421 45543 49479 45549
rect 49421 45540 49433 45543
rect 48832 45512 49433 45540
rect 48832 45500 48838 45512
rect 49421 45509 49433 45512
rect 49467 45509 49479 45543
rect 49421 45503 49479 45509
rect 49602 45500 49608 45552
rect 49660 45540 49666 45552
rect 53193 45543 53251 45549
rect 53193 45540 53205 45543
rect 49660 45512 53205 45540
rect 49660 45500 49666 45512
rect 53193 45509 53205 45512
rect 53239 45540 53251 45543
rect 55769 45543 55827 45549
rect 55769 45540 55781 45543
rect 53239 45512 55781 45540
rect 53239 45509 53251 45512
rect 53193 45503 53251 45509
rect 55769 45509 55781 45512
rect 55815 45509 55827 45543
rect 55769 45503 55827 45509
rect 42981 45475 43039 45481
rect 42981 45441 42993 45475
rect 43027 45441 43039 45475
rect 45922 45472 45928 45484
rect 45883 45444 45928 45472
rect 42981 45435 43039 45441
rect 45922 45432 45928 45444
rect 45980 45432 45986 45484
rect 46017 45475 46075 45481
rect 46017 45441 46029 45475
rect 46063 45472 46075 45475
rect 46474 45472 46480 45484
rect 46063 45444 46480 45472
rect 46063 45441 46075 45444
rect 46017 45435 46075 45441
rect 46474 45432 46480 45444
rect 46532 45432 46538 45484
rect 46753 45475 46811 45481
rect 46753 45441 46765 45475
rect 46799 45472 46811 45475
rect 47118 45472 47124 45484
rect 46799 45444 47124 45472
rect 46799 45441 46811 45444
rect 46753 45435 46811 45441
rect 47118 45432 47124 45444
rect 47176 45432 47182 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 47228 45444 47593 45472
rect 41932 45376 42656 45404
rect 42797 45407 42855 45413
rect 41932 45364 41938 45376
rect 42797 45373 42809 45407
rect 42843 45404 42855 45407
rect 43070 45404 43076 45416
rect 42843 45376 43076 45404
rect 42843 45373 42855 45376
rect 42797 45367 42855 45373
rect 43070 45364 43076 45376
rect 43128 45364 43134 45416
rect 46842 45364 46848 45416
rect 46900 45404 46906 45416
rect 47228 45404 47256 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 47762 45432 47768 45484
rect 47820 45472 47826 45484
rect 47857 45475 47915 45481
rect 47857 45472 47869 45475
rect 47820 45444 47869 45472
rect 47820 45432 47826 45444
rect 47857 45441 47869 45444
rect 47903 45441 47915 45475
rect 47857 45435 47915 45441
rect 48222 45432 48228 45484
rect 48280 45472 48286 45484
rect 48593 45475 48651 45481
rect 48593 45472 48605 45475
rect 48280 45444 48605 45472
rect 48280 45432 48286 45444
rect 48593 45441 48605 45444
rect 48639 45441 48651 45475
rect 48958 45472 48964 45484
rect 48919 45444 48964 45472
rect 48593 45435 48651 45441
rect 48958 45432 48964 45444
rect 49016 45432 49022 45484
rect 49145 45475 49203 45481
rect 49145 45441 49157 45475
rect 49191 45472 49203 45475
rect 49694 45472 49700 45484
rect 49191 45444 49700 45472
rect 49191 45441 49203 45444
rect 49145 45435 49203 45441
rect 49694 45432 49700 45444
rect 49752 45432 49758 45484
rect 51442 45472 51448 45484
rect 51403 45444 51448 45472
rect 51442 45432 51448 45444
rect 51500 45432 51506 45484
rect 55858 45432 55864 45484
rect 55916 45472 55922 45484
rect 55953 45475 56011 45481
rect 55953 45472 55965 45475
rect 55916 45444 55965 45472
rect 55916 45432 55922 45444
rect 55953 45441 55965 45444
rect 55999 45441 56011 45475
rect 55953 45435 56011 45441
rect 56042 45432 56048 45484
rect 56100 45472 56106 45484
rect 56100 45444 56145 45472
rect 56100 45432 56106 45444
rect 47670 45404 47676 45416
rect 46900 45376 47256 45404
rect 47631 45376 47676 45404
rect 46900 45364 46906 45376
rect 47670 45364 47676 45376
rect 47728 45364 47734 45416
rect 48130 45364 48136 45416
rect 48188 45404 48194 45416
rect 51350 45404 51356 45416
rect 48188 45376 51356 45404
rect 48188 45364 48194 45376
rect 51350 45364 51356 45376
rect 51408 45364 51414 45416
rect 51537 45407 51595 45413
rect 51537 45373 51549 45407
rect 51583 45373 51595 45407
rect 51810 45404 51816 45416
rect 51771 45376 51816 45404
rect 51537 45367 51595 45373
rect 43165 45339 43223 45345
rect 43165 45336 43177 45339
rect 40880 45308 43177 45336
rect 43165 45305 43177 45308
rect 43211 45305 43223 45339
rect 43165 45299 43223 45305
rect 47210 45296 47216 45348
rect 47268 45336 47274 45348
rect 48222 45336 48228 45348
rect 47268 45308 48228 45336
rect 47268 45296 47274 45308
rect 48222 45296 48228 45308
rect 48280 45296 48286 45348
rect 49050 45336 49056 45348
rect 49011 45308 49056 45336
rect 49050 45296 49056 45308
rect 49108 45296 49114 45348
rect 51552 45336 51580 45367
rect 51810 45364 51816 45376
rect 51868 45364 51874 45416
rect 51994 45336 52000 45348
rect 51552 45308 52000 45336
rect 51994 45296 52000 45308
rect 52052 45296 52058 45348
rect 41325 45271 41383 45277
rect 41325 45268 41337 45271
rect 38764 45240 41337 45268
rect 41325 45237 41337 45240
rect 41371 45237 41383 45271
rect 41325 45231 41383 45237
rect 42426 45228 42432 45280
rect 42484 45268 42490 45280
rect 45370 45268 45376 45280
rect 42484 45240 45376 45268
rect 42484 45228 42490 45240
rect 45370 45228 45376 45240
rect 45428 45228 45434 45280
rect 45738 45268 45744 45280
rect 45699 45240 45744 45268
rect 45738 45228 45744 45240
rect 45796 45228 45802 45280
rect 46845 45271 46903 45277
rect 46845 45237 46857 45271
rect 46891 45268 46903 45271
rect 47486 45268 47492 45280
rect 46891 45240 47492 45268
rect 46891 45237 46903 45240
rect 46845 45231 46903 45237
rect 47486 45228 47492 45240
rect 47544 45228 47550 45280
rect 47578 45228 47584 45280
rect 47636 45268 47642 45280
rect 47636 45240 47681 45268
rect 47636 45228 47642 45240
rect 52730 45228 52736 45280
rect 52788 45268 52794 45280
rect 53285 45271 53343 45277
rect 53285 45268 53297 45271
rect 52788 45240 53297 45268
rect 52788 45228 52794 45240
rect 53285 45237 53297 45240
rect 53331 45237 53343 45271
rect 53285 45231 53343 45237
rect 55769 45271 55827 45277
rect 55769 45237 55781 45271
rect 55815 45268 55827 45271
rect 55858 45268 55864 45280
rect 55815 45240 55864 45268
rect 55815 45237 55827 45240
rect 55769 45231 55827 45237
rect 55858 45228 55864 45240
rect 55916 45228 55922 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 19245 45067 19303 45073
rect 19245 45033 19257 45067
rect 19291 45064 19303 45067
rect 19334 45064 19340 45076
rect 19291 45036 19340 45064
rect 19291 45033 19303 45036
rect 19245 45027 19303 45033
rect 19334 45024 19340 45036
rect 19392 45024 19398 45076
rect 20162 45064 20168 45076
rect 20123 45036 20168 45064
rect 20162 45024 20168 45036
rect 20220 45024 20226 45076
rect 20533 45067 20591 45073
rect 20533 45033 20545 45067
rect 20579 45064 20591 45067
rect 20622 45064 20628 45076
rect 20579 45036 20628 45064
rect 20579 45033 20591 45036
rect 20533 45027 20591 45033
rect 20622 45024 20628 45036
rect 20680 45024 20686 45076
rect 24854 45024 24860 45076
rect 24912 45064 24918 45076
rect 24949 45067 25007 45073
rect 24949 45064 24961 45067
rect 24912 45036 24961 45064
rect 24912 45024 24918 45036
rect 24949 45033 24961 45036
rect 24995 45064 25007 45067
rect 26050 45064 26056 45076
rect 24995 45036 26056 45064
rect 24995 45033 25007 45036
rect 24949 45027 25007 45033
rect 26050 45024 26056 45036
rect 26108 45024 26114 45076
rect 27341 45067 27399 45073
rect 27341 45033 27353 45067
rect 27387 45064 27399 45067
rect 27706 45064 27712 45076
rect 27387 45036 27712 45064
rect 27387 45033 27399 45036
rect 27341 45027 27399 45033
rect 27706 45024 27712 45036
rect 27764 45024 27770 45076
rect 31018 45064 31024 45076
rect 30760 45036 31024 45064
rect 3418 44956 3424 45008
rect 3476 44996 3482 45008
rect 28994 44996 29000 45008
rect 3476 44968 29000 44996
rect 3476 44956 3482 44968
rect 28994 44956 29000 44968
rect 29052 44996 29058 45008
rect 29270 44996 29276 45008
rect 29052 44968 29276 44996
rect 29052 44956 29058 44968
rect 29270 44956 29276 44968
rect 29328 44956 29334 45008
rect 20257 44931 20315 44937
rect 20257 44897 20269 44931
rect 20303 44928 20315 44931
rect 20438 44928 20444 44940
rect 20303 44900 20444 44928
rect 20303 44897 20315 44900
rect 20257 44891 20315 44897
rect 20438 44888 20444 44900
rect 20496 44888 20502 44940
rect 30760 44937 30788 45036
rect 31018 45024 31024 45036
rect 31076 45024 31082 45076
rect 35434 45024 35440 45076
rect 35492 45064 35498 45076
rect 35492 45036 37136 45064
rect 35492 45024 35498 45036
rect 37108 45005 37136 45036
rect 37182 45024 37188 45076
rect 37240 45064 37246 45076
rect 38010 45064 38016 45076
rect 37240 45036 38016 45064
rect 37240 45024 37246 45036
rect 38010 45024 38016 45036
rect 38068 45024 38074 45076
rect 38378 45064 38384 45076
rect 38339 45036 38384 45064
rect 38378 45024 38384 45036
rect 38436 45024 38442 45076
rect 39114 45064 39120 45076
rect 39075 45036 39120 45064
rect 39114 45024 39120 45036
rect 39172 45024 39178 45076
rect 40313 45067 40371 45073
rect 40313 45033 40325 45067
rect 40359 45064 40371 45067
rect 40954 45064 40960 45076
rect 40359 45036 40960 45064
rect 40359 45033 40371 45036
rect 40313 45027 40371 45033
rect 40954 45024 40960 45036
rect 41012 45024 41018 45076
rect 41322 45024 41328 45076
rect 41380 45064 41386 45076
rect 43438 45064 43444 45076
rect 41380 45036 43444 45064
rect 41380 45024 41386 45036
rect 43438 45024 43444 45036
rect 43496 45024 43502 45076
rect 46566 45064 46572 45076
rect 46527 45036 46572 45064
rect 46566 45024 46572 45036
rect 46624 45024 46630 45076
rect 46937 45067 46995 45073
rect 46937 45033 46949 45067
rect 46983 45064 46995 45067
rect 47118 45064 47124 45076
rect 46983 45036 47124 45064
rect 46983 45033 46995 45036
rect 46937 45027 46995 45033
rect 47118 45024 47124 45036
rect 47176 45024 47182 45076
rect 47670 45024 47676 45076
rect 47728 45064 47734 45076
rect 48133 45067 48191 45073
rect 48133 45064 48145 45067
rect 47728 45036 48145 45064
rect 47728 45024 47734 45036
rect 48133 45033 48145 45036
rect 48179 45033 48191 45067
rect 48133 45027 48191 45033
rect 48222 45024 48228 45076
rect 48280 45064 48286 45076
rect 49510 45064 49516 45076
rect 48280 45036 49516 45064
rect 48280 45024 48286 45036
rect 49510 45024 49516 45036
rect 49568 45024 49574 45076
rect 49605 45067 49663 45073
rect 49605 45033 49617 45067
rect 49651 45064 49663 45067
rect 49694 45064 49700 45076
rect 49651 45036 49700 45064
rect 49651 45033 49663 45036
rect 49605 45027 49663 45033
rect 49694 45024 49700 45036
rect 49752 45064 49758 45076
rect 50706 45064 50712 45076
rect 49752 45036 50712 45064
rect 49752 45024 49758 45036
rect 50706 45024 50712 45036
rect 50764 45024 50770 45076
rect 51350 45024 51356 45076
rect 51408 45064 51414 45076
rect 53469 45067 53527 45073
rect 53469 45064 53481 45067
rect 51408 45036 53481 45064
rect 51408 45024 51414 45036
rect 53469 45033 53481 45036
rect 53515 45033 53527 45067
rect 53469 45027 53527 45033
rect 37093 44999 37151 45005
rect 37093 44965 37105 44999
rect 37139 44965 37151 44999
rect 38657 44999 38715 45005
rect 38657 44996 38669 44999
rect 37093 44959 37151 44965
rect 37292 44968 38669 44996
rect 25869 44931 25927 44937
rect 25869 44928 25881 44931
rect 25056 44900 25881 44928
rect 25056 44872 25084 44900
rect 25869 44897 25881 44900
rect 25915 44897 25927 44931
rect 29917 44931 29975 44937
rect 29917 44928 29929 44931
rect 25869 44891 25927 44897
rect 27540 44900 29929 44928
rect 19426 44860 19432 44872
rect 19387 44832 19432 44860
rect 19426 44820 19432 44832
rect 19484 44820 19490 44872
rect 20349 44863 20407 44869
rect 20349 44829 20361 44863
rect 20395 44860 20407 44863
rect 20530 44860 20536 44872
rect 20395 44832 20536 44860
rect 20395 44829 20407 44832
rect 20349 44823 20407 44829
rect 20530 44820 20536 44832
rect 20588 44820 20594 44872
rect 24670 44860 24676 44872
rect 24631 44832 24676 44860
rect 24670 44820 24676 44832
rect 24728 44820 24734 44872
rect 24762 44820 24768 44872
rect 24820 44860 24826 44872
rect 25038 44860 25044 44872
rect 24820 44832 24865 44860
rect 24951 44832 25044 44860
rect 24820 44820 24826 44832
rect 25038 44820 25044 44832
rect 25096 44820 25102 44872
rect 25590 44860 25596 44872
rect 25551 44832 25596 44860
rect 25590 44820 25596 44832
rect 25648 44820 25654 44872
rect 25682 44820 25688 44872
rect 25740 44860 25746 44872
rect 27540 44869 27568 44900
rect 29917 44897 29929 44900
rect 29963 44897 29975 44931
rect 29917 44891 29975 44897
rect 30745 44931 30803 44937
rect 30745 44897 30757 44931
rect 30791 44897 30803 44931
rect 30745 44891 30803 44897
rect 32030 44888 32036 44940
rect 32088 44928 32094 44940
rect 34606 44928 34612 44940
rect 32088 44900 34612 44928
rect 32088 44888 32094 44900
rect 27525 44863 27583 44869
rect 25740 44832 25785 44860
rect 25740 44820 25746 44832
rect 27525 44829 27537 44863
rect 27571 44829 27583 44863
rect 27525 44823 27583 44829
rect 28169 44863 28227 44869
rect 28169 44829 28181 44863
rect 28215 44860 28227 44863
rect 28258 44860 28264 44872
rect 28215 44832 28264 44860
rect 28215 44829 28227 44832
rect 28169 44823 28227 44829
rect 28258 44820 28264 44832
rect 28316 44820 28322 44872
rect 29086 44820 29092 44872
rect 29144 44860 29150 44872
rect 29549 44863 29607 44869
rect 29549 44860 29561 44863
rect 29144 44832 29561 44860
rect 29144 44820 29150 44832
rect 29549 44829 29561 44832
rect 29595 44829 29607 44863
rect 29549 44823 29607 44829
rect 29733 44863 29791 44869
rect 29733 44829 29745 44863
rect 29779 44860 29791 44863
rect 30282 44860 30288 44872
rect 29779 44832 30288 44860
rect 29779 44829 29791 44832
rect 29733 44823 29791 44829
rect 30282 44820 30288 44832
rect 30340 44820 30346 44872
rect 32214 44860 32220 44872
rect 30392 44832 32220 44860
rect 20073 44795 20131 44801
rect 20073 44761 20085 44795
rect 20119 44792 20131 44795
rect 20254 44792 20260 44804
rect 20119 44764 20260 44792
rect 20119 44761 20131 44764
rect 20073 44755 20131 44761
rect 20254 44752 20260 44764
rect 20312 44752 20318 44804
rect 28810 44792 28816 44804
rect 28771 44764 28816 44792
rect 28810 44752 28816 44764
rect 28868 44792 28874 44804
rect 30392 44792 30420 44832
rect 32214 44820 32220 44832
rect 32272 44820 32278 44872
rect 32398 44820 32404 44872
rect 32456 44860 32462 44872
rect 32815 44863 32873 44869
rect 32815 44860 32827 44863
rect 32456 44832 32827 44860
rect 32456 44820 32462 44832
rect 32815 44829 32827 44832
rect 32861 44829 32873 44863
rect 32950 44860 32956 44872
rect 32911 44832 32956 44860
rect 32815 44823 32873 44829
rect 32950 44820 32956 44832
rect 33008 44820 33014 44872
rect 33060 44869 33088 44900
rect 34606 44888 34612 44900
rect 34664 44888 34670 44940
rect 37292 44937 37320 44968
rect 38657 44965 38669 44968
rect 38703 44965 38715 44999
rect 38657 44959 38715 44965
rect 41598 44956 41604 45008
rect 41656 44996 41662 45008
rect 49418 44996 49424 45008
rect 41656 44968 49424 44996
rect 41656 44956 41662 44968
rect 49418 44956 49424 44968
rect 49476 44956 49482 45008
rect 55490 44996 55496 45008
rect 55451 44968 55496 44996
rect 55490 44956 55496 44968
rect 55548 44956 55554 45008
rect 57790 44996 57796 45008
rect 56336 44968 57796 44996
rect 37277 44931 37335 44937
rect 37277 44897 37289 44931
rect 37323 44897 37335 44931
rect 37277 44891 37335 44897
rect 37369 44931 37427 44937
rect 37369 44897 37381 44931
rect 37415 44928 37427 44931
rect 37734 44928 37740 44940
rect 37415 44900 37740 44928
rect 37415 44897 37427 44900
rect 37369 44891 37427 44897
rect 37734 44888 37740 44900
rect 37792 44888 37798 44940
rect 37918 44888 37924 44940
rect 37976 44928 37982 44940
rect 37976 44900 39436 44928
rect 37976 44888 37982 44900
rect 33045 44863 33103 44869
rect 33045 44829 33057 44863
rect 33091 44829 33103 44863
rect 33045 44823 33103 44829
rect 33229 44863 33287 44869
rect 33229 44829 33241 44863
rect 33275 44829 33287 44863
rect 33229 44823 33287 44829
rect 28868 44764 30420 44792
rect 31012 44795 31070 44801
rect 28868 44752 28874 44764
rect 31012 44761 31024 44795
rect 31058 44792 31070 44795
rect 32585 44795 32643 44801
rect 32585 44792 32597 44795
rect 31058 44764 32597 44792
rect 31058 44761 31070 44764
rect 31012 44755 31070 44761
rect 32585 44761 32597 44764
rect 32631 44761 32643 44795
rect 33244 44792 33272 44823
rect 33502 44820 33508 44872
rect 33560 44860 33566 44872
rect 34701 44863 34759 44869
rect 34701 44860 34713 44863
rect 33560 44832 34713 44860
rect 33560 44820 33566 44832
rect 34701 44829 34713 44832
rect 34747 44829 34759 44863
rect 34701 44823 34759 44829
rect 34968 44863 35026 44869
rect 34968 44829 34980 44863
rect 35014 44860 35026 44863
rect 35710 44860 35716 44872
rect 35014 44832 35716 44860
rect 35014 44829 35026 44832
rect 34968 44823 35026 44829
rect 35710 44820 35716 44832
rect 35768 44820 35774 44872
rect 37461 44863 37519 44869
rect 37461 44829 37473 44863
rect 37507 44829 37519 44863
rect 37461 44823 37519 44829
rect 37476 44792 37504 44823
rect 37550 44820 37556 44872
rect 37608 44860 37614 44872
rect 37608 44832 37653 44860
rect 37608 44820 37614 44832
rect 37826 44820 37832 44872
rect 37884 44860 37890 44872
rect 38105 44863 38163 44869
rect 38105 44860 38117 44863
rect 37884 44832 38117 44860
rect 37884 44820 37890 44832
rect 38105 44829 38117 44832
rect 38151 44829 38163 44863
rect 38105 44823 38163 44829
rect 38194 44820 38200 44872
rect 38252 44860 38258 44872
rect 38378 44860 38384 44872
rect 38252 44832 38384 44860
rect 38252 44820 38258 44832
rect 38378 44820 38384 44832
rect 38436 44820 38442 44872
rect 38654 44820 38660 44872
rect 38712 44860 38718 44872
rect 39117 44863 39175 44869
rect 39117 44860 39129 44863
rect 38712 44832 39129 44860
rect 38712 44820 38718 44832
rect 39117 44829 39129 44832
rect 39163 44829 39175 44863
rect 39298 44860 39304 44872
rect 39259 44832 39304 44860
rect 39117 44823 39175 44829
rect 39298 44820 39304 44832
rect 39356 44820 39362 44872
rect 39408 44860 39436 44900
rect 40126 44888 40132 44940
rect 40184 44928 40190 44940
rect 49050 44928 49056 44940
rect 40184 44900 40632 44928
rect 40184 44888 40190 44900
rect 39666 44860 39672 44872
rect 39408 44832 39672 44860
rect 39666 44820 39672 44832
rect 39724 44820 39730 44872
rect 39850 44820 39856 44872
rect 39908 44860 39914 44872
rect 40497 44863 40555 44869
rect 40497 44860 40509 44863
rect 39908 44832 40509 44860
rect 39908 44820 39914 44832
rect 40497 44829 40509 44832
rect 40543 44829 40555 44863
rect 40604 44860 40632 44900
rect 42260 44900 49056 44928
rect 40865 44863 40923 44869
rect 40865 44860 40877 44863
rect 40604 44832 40877 44860
rect 40497 44823 40555 44829
rect 40865 44829 40877 44832
rect 40911 44829 40923 44863
rect 40865 44823 40923 44829
rect 40957 44863 41015 44869
rect 40957 44829 40969 44863
rect 41003 44860 41015 44863
rect 41046 44860 41052 44872
rect 41003 44832 41052 44860
rect 41003 44829 41015 44832
rect 40957 44823 41015 44829
rect 41046 44820 41052 44832
rect 41104 44820 41110 44872
rect 42153 44863 42211 44869
rect 42153 44829 42165 44863
rect 42199 44862 42211 44863
rect 42260 44862 42288 44900
rect 49050 44888 49056 44900
rect 49108 44888 49114 44940
rect 49237 44931 49295 44937
rect 49237 44897 49249 44931
rect 49283 44928 49295 44931
rect 49326 44928 49332 44940
rect 49283 44900 49332 44928
rect 49283 44897 49295 44900
rect 49237 44891 49295 44897
rect 49326 44888 49332 44900
rect 49384 44888 49390 44940
rect 49510 44888 49516 44940
rect 49568 44928 49574 44940
rect 52638 44928 52644 44940
rect 49568 44900 51672 44928
rect 49568 44888 49574 44900
rect 42199 44834 42288 44862
rect 42426 44860 42432 44872
rect 42199 44829 42211 44834
rect 42387 44832 42432 44860
rect 42153 44823 42211 44829
rect 42426 44820 42432 44832
rect 42484 44820 42490 44872
rect 43257 44863 43315 44869
rect 43257 44860 43269 44863
rect 42536 44832 43269 44860
rect 38470 44792 38476 44804
rect 33244 44764 37320 44792
rect 37476 44764 38476 44792
rect 32585 44755 32643 44761
rect 24210 44684 24216 44736
rect 24268 44724 24274 44736
rect 24489 44727 24547 44733
rect 24489 44724 24501 44727
rect 24268 44696 24501 44724
rect 24268 44684 24274 44696
rect 24489 44693 24501 44696
rect 24535 44693 24547 44727
rect 24489 44687 24547 44693
rect 32125 44727 32183 44733
rect 32125 44693 32137 44727
rect 32171 44724 32183 44727
rect 32950 44724 32956 44736
rect 32171 44696 32956 44724
rect 32171 44693 32183 44696
rect 32125 44687 32183 44693
rect 32950 44684 32956 44696
rect 33008 44684 33014 44736
rect 34330 44684 34336 44736
rect 34388 44724 34394 44736
rect 35618 44724 35624 44736
rect 34388 44696 35624 44724
rect 34388 44684 34394 44696
rect 35618 44684 35624 44696
rect 35676 44724 35682 44736
rect 36081 44727 36139 44733
rect 36081 44724 36093 44727
rect 35676 44696 36093 44724
rect 35676 44684 35682 44696
rect 36081 44693 36093 44696
rect 36127 44693 36139 44727
rect 37292 44724 37320 44764
rect 38470 44752 38476 44764
rect 38528 44752 38534 44804
rect 40586 44792 40592 44804
rect 40547 44764 40592 44792
rect 40586 44752 40592 44764
rect 40644 44752 40650 44804
rect 40681 44795 40739 44801
rect 40681 44761 40693 44795
rect 40727 44792 40739 44795
rect 42242 44792 42248 44804
rect 40727 44764 42248 44792
rect 40727 44761 40739 44764
rect 40681 44755 40739 44761
rect 42242 44752 42248 44764
rect 42300 44792 42306 44804
rect 42536 44792 42564 44832
rect 43257 44829 43269 44832
rect 43303 44829 43315 44863
rect 43257 44823 43315 44829
rect 44082 44820 44088 44872
rect 44140 44860 44146 44872
rect 45465 44863 45523 44869
rect 45465 44860 45477 44863
rect 44140 44832 45477 44860
rect 44140 44820 44146 44832
rect 45465 44829 45477 44832
rect 45511 44829 45523 44863
rect 46474 44860 46480 44872
rect 46435 44832 46480 44860
rect 45465 44823 45523 44829
rect 46474 44820 46480 44832
rect 46532 44820 46538 44872
rect 47026 44820 47032 44872
rect 47084 44860 47090 44872
rect 47765 44863 47823 44869
rect 47765 44860 47777 44863
rect 47084 44832 47777 44860
rect 47084 44820 47090 44832
rect 47765 44829 47777 44832
rect 47811 44829 47823 44863
rect 47765 44823 47823 44829
rect 47949 44863 48007 44869
rect 47949 44829 47961 44863
rect 47995 44860 48007 44863
rect 48222 44860 48228 44872
rect 47995 44832 48228 44860
rect 47995 44829 48007 44832
rect 47949 44823 48007 44829
rect 48222 44820 48228 44832
rect 48280 44820 48286 44872
rect 49418 44860 49424 44872
rect 49379 44832 49424 44860
rect 49418 44820 49424 44832
rect 49476 44820 49482 44872
rect 51644 44869 51672 44900
rect 51920 44900 52644 44928
rect 51920 44869 51948 44900
rect 52638 44888 52644 44900
rect 52696 44888 52702 44940
rect 53834 44928 53840 44940
rect 53024 44900 53840 44928
rect 50709 44863 50767 44869
rect 50709 44829 50721 44863
rect 50755 44829 50767 44863
rect 50709 44823 50767 44829
rect 50985 44863 51043 44869
rect 50985 44829 50997 44863
rect 51031 44860 51043 44863
rect 51445 44863 51503 44869
rect 51445 44860 51457 44863
rect 51031 44832 51457 44860
rect 51031 44829 51043 44832
rect 50985 44823 51043 44829
rect 51445 44829 51457 44832
rect 51491 44829 51503 44863
rect 51445 44823 51503 44829
rect 51629 44863 51687 44869
rect 51629 44829 51641 44863
rect 51675 44829 51687 44863
rect 51629 44823 51687 44829
rect 51905 44863 51963 44869
rect 51905 44829 51917 44863
rect 51951 44829 51963 44863
rect 52086 44860 52092 44872
rect 52047 44832 52092 44860
rect 51905 44823 51963 44829
rect 42886 44792 42892 44804
rect 42300 44764 42564 44792
rect 42847 44764 42892 44792
rect 42300 44752 42306 44764
rect 42886 44752 42892 44764
rect 42944 44752 42950 44804
rect 42978 44752 42984 44804
rect 43036 44792 43042 44804
rect 43073 44795 43131 44801
rect 43073 44792 43085 44795
rect 43036 44764 43085 44792
rect 43036 44752 43042 44764
rect 43073 44761 43085 44764
rect 43119 44761 43131 44795
rect 43073 44755 43131 44761
rect 43162 44752 43168 44804
rect 43220 44792 43226 44804
rect 44100 44792 44128 44820
rect 43220 44764 44128 44792
rect 43220 44752 43226 44764
rect 44174 44752 44180 44804
rect 44232 44792 44238 44804
rect 50724 44792 50752 44823
rect 44232 44764 50752 44792
rect 51644 44792 51672 44823
rect 52086 44820 52092 44832
rect 52144 44820 52150 44872
rect 52730 44860 52736 44872
rect 52196 44832 52736 44860
rect 52196 44792 52224 44832
rect 52730 44820 52736 44832
rect 52788 44820 52794 44872
rect 53024 44869 53052 44900
rect 53834 44888 53840 44900
rect 53892 44888 53898 44940
rect 56042 44928 56048 44940
rect 55508 44900 56048 44928
rect 53009 44863 53067 44869
rect 53009 44829 53021 44863
rect 53055 44829 53067 44863
rect 53009 44823 53067 44829
rect 53469 44863 53527 44869
rect 53469 44829 53481 44863
rect 53515 44829 53527 44863
rect 53650 44860 53656 44872
rect 53611 44832 53656 44860
rect 53469 44823 53527 44829
rect 51644 44764 52224 44792
rect 52549 44795 52607 44801
rect 44232 44752 44238 44764
rect 52549 44761 52561 44795
rect 52595 44792 52607 44795
rect 53484 44792 53512 44823
rect 53650 44820 53656 44832
rect 53708 44820 53714 44872
rect 55508 44869 55536 44900
rect 56042 44888 56048 44900
rect 56100 44888 56106 44940
rect 56336 44937 56364 44968
rect 57790 44956 57796 44968
rect 57848 44956 57854 45008
rect 56321 44931 56379 44937
rect 56321 44897 56333 44931
rect 56367 44897 56379 44931
rect 56321 44891 56379 44897
rect 56505 44931 56563 44937
rect 56505 44897 56517 44931
rect 56551 44928 56563 44931
rect 57054 44928 57060 44940
rect 56551 44900 57060 44928
rect 56551 44897 56563 44900
rect 56505 44891 56563 44897
rect 57054 44888 57060 44900
rect 57112 44888 57118 44940
rect 57882 44928 57888 44940
rect 57843 44900 57888 44928
rect 57882 44888 57888 44900
rect 57940 44888 57946 44940
rect 55493 44863 55551 44869
rect 55493 44829 55505 44863
rect 55539 44829 55551 44863
rect 55493 44823 55551 44829
rect 55677 44863 55735 44869
rect 55677 44829 55689 44863
rect 55723 44829 55735 44863
rect 55858 44860 55864 44872
rect 55819 44832 55864 44860
rect 55677 44823 55735 44829
rect 52595 44764 53512 44792
rect 55692 44792 55720 44823
rect 55858 44820 55864 44832
rect 55916 44820 55922 44872
rect 55766 44792 55772 44804
rect 55692 44764 55772 44792
rect 52595 44761 52607 44764
rect 52549 44755 52607 44761
rect 55766 44752 55772 44764
rect 55824 44752 55830 44804
rect 41969 44727 42027 44733
rect 41969 44724 41981 44727
rect 37292 44696 41981 44724
rect 36081 44687 36139 44693
rect 41969 44693 41981 44696
rect 42015 44693 42027 44727
rect 42334 44724 42340 44736
rect 42295 44696 42340 44724
rect 41969 44687 42027 44693
rect 42334 44684 42340 44696
rect 42392 44684 42398 44736
rect 42518 44684 42524 44736
rect 42576 44724 42582 44736
rect 44358 44724 44364 44736
rect 42576 44696 44364 44724
rect 42576 44684 42582 44696
rect 44358 44684 44364 44696
rect 44416 44684 44422 44736
rect 45554 44724 45560 44736
rect 45515 44696 45560 44724
rect 45554 44684 45560 44696
rect 45612 44684 45618 44736
rect 49694 44684 49700 44736
rect 49752 44724 49758 44736
rect 50525 44727 50583 44733
rect 50525 44724 50537 44727
rect 49752 44696 50537 44724
rect 49752 44684 49758 44696
rect 50525 44693 50537 44696
rect 50571 44693 50583 44727
rect 50890 44724 50896 44736
rect 50851 44696 50896 44724
rect 50525 44687 50583 44693
rect 50890 44684 50896 44696
rect 50948 44684 50954 44736
rect 52914 44724 52920 44736
rect 52875 44696 52920 44724
rect 52914 44684 52920 44696
rect 52972 44684 52978 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 19521 44523 19579 44529
rect 19521 44489 19533 44523
rect 19567 44520 19579 44523
rect 19978 44520 19984 44532
rect 19567 44492 19984 44520
rect 19567 44489 19579 44492
rect 19521 44483 19579 44489
rect 19978 44480 19984 44492
rect 20036 44480 20042 44532
rect 24762 44480 24768 44532
rect 24820 44480 24826 44532
rect 38562 44480 38568 44532
rect 38620 44520 38626 44532
rect 39685 44523 39743 44529
rect 39685 44520 39697 44523
rect 38620 44492 39697 44520
rect 38620 44480 38626 44492
rect 39685 44489 39697 44492
rect 39731 44489 39743 44523
rect 39850 44520 39856 44532
rect 39811 44492 39856 44520
rect 39685 44483 39743 44489
rect 39850 44480 39856 44492
rect 39908 44480 39914 44532
rect 40862 44480 40868 44532
rect 40920 44520 40926 44532
rect 41782 44520 41788 44532
rect 40920 44492 41788 44520
rect 40920 44480 40926 44492
rect 41782 44480 41788 44492
rect 41840 44480 41846 44532
rect 42978 44520 42984 44532
rect 42644 44492 42984 44520
rect 2038 44412 2044 44464
rect 2096 44452 2102 44464
rect 2682 44452 2688 44464
rect 2096 44424 2688 44452
rect 2096 44412 2102 44424
rect 2682 44412 2688 44424
rect 2740 44412 2746 44464
rect 24780 44452 24808 44480
rect 24688 44424 24808 44452
rect 19705 44387 19763 44393
rect 19705 44353 19717 44387
rect 19751 44384 19763 44387
rect 20070 44384 20076 44396
rect 19751 44356 20076 44384
rect 19751 44353 19763 44356
rect 19705 44347 19763 44353
rect 20070 44344 20076 44356
rect 20128 44344 20134 44396
rect 24688 44393 24716 44424
rect 27614 44412 27620 44464
rect 27672 44452 27678 44464
rect 31018 44452 31024 44464
rect 27672 44424 31024 44452
rect 27672 44412 27678 44424
rect 24673 44387 24731 44393
rect 24673 44353 24685 44387
rect 24719 44353 24731 44387
rect 24673 44347 24731 44353
rect 24765 44387 24823 44393
rect 24765 44353 24777 44387
rect 24811 44384 24823 44387
rect 24854 44384 24860 44396
rect 24811 44356 24860 44384
rect 24811 44353 24823 44356
rect 24765 44347 24823 44353
rect 24854 44344 24860 44356
rect 24912 44344 24918 44396
rect 25038 44384 25044 44396
rect 24999 44356 25044 44384
rect 25038 44344 25044 44356
rect 25096 44344 25102 44396
rect 28092 44393 28120 44424
rect 31018 44412 31024 44424
rect 31076 44412 31082 44464
rect 32030 44412 32036 44464
rect 32088 44452 32094 44464
rect 33772 44455 33830 44461
rect 32088 44424 32628 44452
rect 32088 44412 32094 44424
rect 28077 44387 28135 44393
rect 28077 44353 28089 44387
rect 28123 44353 28135 44387
rect 28077 44347 28135 44353
rect 28344 44387 28402 44393
rect 28344 44353 28356 44387
rect 28390 44384 28402 44387
rect 29454 44384 29460 44396
rect 28390 44356 29460 44384
rect 28390 44353 28402 44356
rect 28344 44347 28402 44353
rect 29454 44344 29460 44356
rect 29512 44344 29518 44396
rect 32398 44384 32404 44396
rect 32359 44356 32404 44384
rect 32398 44344 32404 44356
rect 32456 44344 32462 44396
rect 32600 44393 32628 44424
rect 33772 44421 33784 44455
rect 33818 44452 33830 44455
rect 35345 44455 35403 44461
rect 35345 44452 35357 44455
rect 33818 44424 35357 44452
rect 33818 44421 33830 44424
rect 33772 44415 33830 44421
rect 35345 44421 35357 44424
rect 35391 44421 35403 44455
rect 35345 44415 35403 44421
rect 37826 44412 37832 44464
rect 37884 44452 37890 44464
rect 39114 44452 39120 44464
rect 37884 44424 39120 44452
rect 37884 44412 37890 44424
rect 39114 44412 39120 44424
rect 39172 44452 39178 44464
rect 39485 44455 39543 44461
rect 39485 44452 39497 44455
rect 39172 44424 39497 44452
rect 39172 44412 39178 44424
rect 39485 44421 39497 44424
rect 39531 44421 39543 44455
rect 39485 44415 39543 44421
rect 40586 44412 40592 44464
rect 40644 44452 40650 44464
rect 41417 44455 41475 44461
rect 41417 44452 41429 44455
rect 40644 44424 41429 44452
rect 40644 44412 40650 44424
rect 41417 44421 41429 44424
rect 41463 44421 41475 44455
rect 41417 44415 41475 44421
rect 32493 44387 32551 44393
rect 32493 44353 32505 44387
rect 32539 44353 32551 44387
rect 32493 44347 32551 44353
rect 32585 44387 32643 44393
rect 32585 44353 32597 44387
rect 32631 44353 32643 44387
rect 32766 44384 32772 44396
rect 32727 44356 32772 44384
rect 32585 44347 32643 44353
rect 32508 44316 32536 44347
rect 32766 44344 32772 44356
rect 32824 44344 32830 44396
rect 33502 44384 33508 44396
rect 33463 44356 33508 44384
rect 33502 44344 33508 44356
rect 33560 44344 33566 44396
rect 35526 44344 35532 44396
rect 35584 44384 35590 44396
rect 35621 44387 35679 44393
rect 35621 44384 35633 44387
rect 35584 44356 35633 44384
rect 35584 44344 35590 44356
rect 35621 44353 35633 44356
rect 35667 44353 35679 44387
rect 35621 44347 35679 44353
rect 35713 44387 35771 44393
rect 35713 44353 35725 44387
rect 35759 44353 35771 44387
rect 35713 44347 35771 44353
rect 35728 44316 35756 44347
rect 35802 44344 35808 44396
rect 35860 44384 35866 44396
rect 35986 44384 35992 44396
rect 35860 44356 35905 44384
rect 35947 44356 35992 44384
rect 35860 44344 35866 44356
rect 35986 44344 35992 44356
rect 36044 44344 36050 44396
rect 39298 44344 39304 44396
rect 39356 44384 39362 44396
rect 41138 44384 41144 44396
rect 39356 44356 41144 44384
rect 39356 44344 39362 44356
rect 41138 44344 41144 44356
rect 41196 44344 41202 44396
rect 41322 44384 41328 44396
rect 41283 44356 41328 44384
rect 41322 44344 41328 44356
rect 41380 44384 41386 44396
rect 41874 44384 41880 44396
rect 41380 44356 41880 44384
rect 41380 44344 41386 44356
rect 41874 44344 41880 44356
rect 41932 44344 41938 44396
rect 42644 44393 42672 44492
rect 42978 44480 42984 44492
rect 43036 44520 43042 44532
rect 43438 44520 43444 44532
rect 43036 44492 43444 44520
rect 43036 44480 43042 44492
rect 43438 44480 43444 44492
rect 43496 44480 43502 44532
rect 43717 44523 43775 44529
rect 43717 44489 43729 44523
rect 43763 44520 43775 44523
rect 44174 44520 44180 44532
rect 43763 44492 44180 44520
rect 43763 44489 43775 44492
rect 43717 44483 43775 44489
rect 44174 44480 44180 44492
rect 44232 44480 44238 44532
rect 47854 44520 47860 44532
rect 45572 44492 47860 44520
rect 44358 44412 44364 44464
rect 44416 44452 44422 44464
rect 45572 44461 45600 44492
rect 47854 44480 47860 44492
rect 47912 44480 47918 44532
rect 48222 44520 48228 44532
rect 48183 44492 48228 44520
rect 48222 44480 48228 44492
rect 48280 44480 48286 44532
rect 48958 44480 48964 44532
rect 49016 44520 49022 44532
rect 49237 44523 49295 44529
rect 49237 44520 49249 44523
rect 49016 44492 49249 44520
rect 49016 44480 49022 44492
rect 49237 44489 49249 44492
rect 49283 44489 49295 44523
rect 49237 44483 49295 44489
rect 50890 44480 50896 44532
rect 50948 44520 50954 44532
rect 52089 44523 52147 44529
rect 52089 44520 52101 44523
rect 50948 44492 52101 44520
rect 50948 44480 50954 44492
rect 52089 44489 52101 44492
rect 52135 44520 52147 44523
rect 52914 44520 52920 44532
rect 52135 44492 52920 44520
rect 52135 44489 52147 44492
rect 52089 44483 52147 44489
rect 52914 44480 52920 44492
rect 52972 44480 52978 44532
rect 53650 44520 53656 44532
rect 53611 44492 53656 44520
rect 53650 44480 53656 44492
rect 53708 44520 53714 44532
rect 53708 44492 54524 44520
rect 53708 44480 53714 44492
rect 45557 44455 45615 44461
rect 45557 44452 45569 44455
rect 44416 44424 45569 44452
rect 44416 44412 44422 44424
rect 45557 44421 45569 44424
rect 45603 44421 45615 44455
rect 47302 44452 47308 44464
rect 45557 44415 45615 44421
rect 45664 44424 47308 44452
rect 42613 44387 42672 44393
rect 42613 44384 42625 44387
rect 42168 44356 42625 44384
rect 32416 44288 32536 44316
rect 34900 44288 35756 44316
rect 32416 44260 32444 44288
rect 24670 44208 24676 44260
rect 24728 44248 24734 44260
rect 24949 44251 25007 44257
rect 24949 44248 24961 44251
rect 24728 44220 24961 44248
rect 24728 44208 24734 44220
rect 24949 44217 24961 44220
rect 24995 44217 25007 44251
rect 24949 44211 25007 44217
rect 32398 44208 32404 44260
rect 32456 44208 32462 44260
rect 2958 44140 2964 44192
rect 3016 44180 3022 44192
rect 3418 44180 3424 44192
rect 3016 44152 3424 44180
rect 3016 44140 3022 44152
rect 3418 44140 3424 44152
rect 3476 44140 3482 44192
rect 24394 44140 24400 44192
rect 24452 44180 24458 44192
rect 24489 44183 24547 44189
rect 24489 44180 24501 44183
rect 24452 44152 24501 44180
rect 24452 44140 24458 44152
rect 24489 44149 24501 44152
rect 24535 44149 24547 44183
rect 24489 44143 24547 44149
rect 29457 44183 29515 44189
rect 29457 44149 29469 44183
rect 29503 44180 29515 44183
rect 30190 44180 30196 44192
rect 29503 44152 30196 44180
rect 29503 44149 29515 44152
rect 29457 44143 29515 44149
rect 30190 44140 30196 44152
rect 30248 44140 30254 44192
rect 32122 44180 32128 44192
rect 32083 44152 32128 44180
rect 32122 44140 32128 44152
rect 32180 44140 32186 44192
rect 34514 44140 34520 44192
rect 34572 44180 34578 44192
rect 34900 44189 34928 44288
rect 38378 44276 38384 44328
rect 38436 44316 38442 44328
rect 42168 44316 42196 44356
rect 42613 44353 42625 44356
rect 42659 44356 42672 44387
rect 42705 44387 42763 44393
rect 42659 44353 42671 44356
rect 42613 44347 42671 44353
rect 42705 44353 42717 44387
rect 42751 44353 42763 44387
rect 42886 44384 42892 44396
rect 42799 44356 42892 44384
rect 42705 44347 42763 44353
rect 38436 44288 42196 44316
rect 38436 44276 38442 44288
rect 42720 44260 42748 44347
rect 42886 44344 42892 44356
rect 42944 44344 42950 44396
rect 42981 44387 43039 44393
rect 42981 44353 42993 44387
rect 43027 44384 43039 44387
rect 43162 44384 43168 44396
rect 43027 44356 43168 44384
rect 43027 44353 43039 44356
rect 42981 44347 43039 44353
rect 43162 44344 43168 44356
rect 43220 44344 43226 44396
rect 43441 44387 43499 44393
rect 43441 44353 43453 44387
rect 43487 44384 43499 44387
rect 43898 44384 43904 44396
rect 43487 44356 43904 44384
rect 43487 44353 43499 44356
rect 43441 44347 43499 44353
rect 43898 44344 43904 44356
rect 43956 44344 43962 44396
rect 44818 44384 44824 44396
rect 44779 44356 44824 44384
rect 44818 44344 44824 44356
rect 44876 44344 44882 44396
rect 45005 44387 45063 44393
rect 45005 44353 45017 44387
rect 45051 44384 45063 44387
rect 45462 44384 45468 44396
rect 45051 44356 45468 44384
rect 45051 44353 45063 44356
rect 45005 44347 45063 44353
rect 45462 44344 45468 44356
rect 45520 44384 45526 44396
rect 45664 44384 45692 44424
rect 45520 44356 45692 44384
rect 46401 44390 46429 44424
rect 47302 44412 47308 44424
rect 47360 44412 47366 44464
rect 49418 44452 49424 44464
rect 49160 44424 49424 44452
rect 46478 44390 46536 44393
rect 46401 44387 46536 44390
rect 46401 44362 46490 44387
rect 45520 44344 45526 44356
rect 46478 44353 46490 44362
rect 46524 44353 46536 44387
rect 46478 44347 46536 44353
rect 46658 44344 46664 44396
rect 46716 44384 46722 44396
rect 47857 44387 47915 44393
rect 46716 44356 46761 44384
rect 46716 44344 46722 44356
rect 47857 44353 47869 44387
rect 47903 44353 47915 44387
rect 47857 44347 47915 44353
rect 48041 44387 48099 44393
rect 48041 44353 48053 44387
rect 48087 44384 48099 44387
rect 48314 44384 48320 44396
rect 48087 44356 48320 44384
rect 48087 44353 48099 44356
rect 48041 44347 48099 44353
rect 42904 44316 42932 44344
rect 43254 44316 43260 44328
rect 42904 44288 43260 44316
rect 43254 44276 43260 44288
rect 43312 44276 43318 44328
rect 43530 44316 43536 44328
rect 43491 44288 43536 44316
rect 43530 44276 43536 44288
rect 43588 44276 43594 44328
rect 43714 44316 43720 44328
rect 43675 44288 43720 44316
rect 43714 44276 43720 44288
rect 43772 44276 43778 44328
rect 46385 44319 46443 44325
rect 46385 44285 46397 44319
rect 46431 44285 46443 44319
rect 46385 44279 46443 44285
rect 38286 44208 38292 44260
rect 38344 44248 38350 44260
rect 41230 44248 41236 44260
rect 38344 44220 41236 44248
rect 38344 44208 38350 44220
rect 41230 44208 41236 44220
rect 41288 44208 41294 44260
rect 41966 44208 41972 44260
rect 42024 44248 42030 44260
rect 42702 44248 42708 44260
rect 42024 44220 42708 44248
rect 42024 44208 42030 44220
rect 42702 44208 42708 44220
rect 42760 44208 42766 44260
rect 45741 44251 45799 44257
rect 45741 44217 45753 44251
rect 45787 44248 45799 44251
rect 45830 44248 45836 44260
rect 45787 44220 45836 44248
rect 45787 44217 45799 44220
rect 45741 44211 45799 44217
rect 45830 44208 45836 44220
rect 45888 44208 45894 44260
rect 46401 44248 46429 44279
rect 46566 44276 46572 44328
rect 46624 44316 46630 44328
rect 47872 44316 47900 44347
rect 48314 44344 48320 44356
rect 48372 44384 48378 44396
rect 48774 44384 48780 44396
rect 48372 44356 48780 44384
rect 48372 44344 48378 44356
rect 48774 44344 48780 44356
rect 48832 44344 48838 44396
rect 49160 44393 49188 44424
rect 49418 44412 49424 44424
rect 49476 44452 49482 44464
rect 50157 44455 50215 44461
rect 50157 44452 50169 44455
rect 49476 44424 50169 44452
rect 49476 44412 49482 44424
rect 50157 44421 50169 44424
rect 50203 44421 50215 44455
rect 50982 44452 50988 44464
rect 50943 44424 50988 44452
rect 50157 44415 50215 44421
rect 50982 44412 50988 44424
rect 51040 44412 51046 44464
rect 51169 44455 51227 44461
rect 51169 44421 51181 44455
rect 51215 44452 51227 44455
rect 51442 44452 51448 44464
rect 51215 44424 51448 44452
rect 51215 44421 51227 44424
rect 51169 44415 51227 44421
rect 51442 44412 51448 44424
rect 51500 44452 51506 44464
rect 52932 44452 52960 44480
rect 54496 44461 54524 44492
rect 54481 44455 54539 44461
rect 51500 44424 52776 44452
rect 52932 44424 53788 44452
rect 51500 44412 51506 44424
rect 49145 44387 49203 44393
rect 49145 44353 49157 44387
rect 49191 44353 49203 44387
rect 49326 44384 49332 44396
rect 49287 44356 49332 44384
rect 49145 44347 49203 44353
rect 49326 44344 49332 44356
rect 49384 44344 49390 44396
rect 50062 44384 50068 44396
rect 50023 44356 50068 44384
rect 50062 44344 50068 44356
rect 50120 44344 50126 44396
rect 50249 44387 50307 44393
rect 50249 44353 50261 44387
rect 50295 44384 50307 44387
rect 50801 44387 50859 44393
rect 50801 44384 50813 44387
rect 50295 44356 50813 44384
rect 50295 44353 50307 44356
rect 50249 44347 50307 44353
rect 50801 44353 50813 44356
rect 50847 44353 50859 44387
rect 50801 44347 50859 44353
rect 51997 44387 52055 44393
rect 51997 44353 52009 44387
rect 52043 44353 52055 44387
rect 51997 44347 52055 44353
rect 48222 44316 48228 44328
rect 46624 44288 46669 44316
rect 47872 44288 48228 44316
rect 46624 44276 46630 44288
rect 48222 44276 48228 44288
rect 48280 44276 48286 44328
rect 50816 44316 50844 44347
rect 50890 44316 50896 44328
rect 50816 44288 50896 44316
rect 50890 44276 50896 44288
rect 50948 44276 50954 44328
rect 52012 44316 52040 44347
rect 52086 44344 52092 44396
rect 52144 44384 52150 44396
rect 52748 44393 52776 44424
rect 53760 44393 53788 44424
rect 54481 44421 54493 44455
rect 54527 44421 54539 44455
rect 54481 44415 54539 44421
rect 54665 44455 54723 44461
rect 54665 44421 54677 44455
rect 54711 44452 54723 44455
rect 55122 44452 55128 44464
rect 54711 44424 55128 44452
rect 54711 44421 54723 44424
rect 54665 44415 54723 44421
rect 52181 44387 52239 44393
rect 52181 44384 52193 44387
rect 52144 44356 52193 44384
rect 52144 44344 52150 44356
rect 52181 44353 52193 44356
rect 52227 44353 52239 44387
rect 52181 44347 52239 44353
rect 52733 44387 52791 44393
rect 52733 44353 52745 44387
rect 52779 44353 52791 44387
rect 52733 44347 52791 44353
rect 52917 44387 52975 44393
rect 52917 44353 52929 44387
rect 52963 44353 52975 44387
rect 52917 44347 52975 44353
rect 53561 44387 53619 44393
rect 53561 44353 53573 44387
rect 53607 44353 53619 44387
rect 53561 44347 53619 44353
rect 53745 44387 53803 44393
rect 53745 44353 53757 44387
rect 53791 44353 53803 44387
rect 53745 44347 53803 44353
rect 52638 44316 52644 44328
rect 52012 44288 52644 44316
rect 52638 44276 52644 44288
rect 52696 44276 52702 44328
rect 47118 44248 47124 44260
rect 46401 44220 47124 44248
rect 47118 44208 47124 44220
rect 47176 44208 47182 44260
rect 52086 44208 52092 44260
rect 52144 44248 52150 44260
rect 52932 44248 52960 44347
rect 53576 44316 53604 44347
rect 53834 44316 53840 44328
rect 53576 44288 53840 44316
rect 53834 44276 53840 44288
rect 53892 44276 53898 44328
rect 54496 44316 54524 44415
rect 55122 44412 55128 44424
rect 55180 44452 55186 44464
rect 55217 44455 55275 44461
rect 55217 44452 55229 44455
rect 55180 44424 55229 44452
rect 55180 44412 55186 44424
rect 55217 44421 55229 44424
rect 55263 44421 55275 44455
rect 55217 44415 55275 44421
rect 55861 44455 55919 44461
rect 55861 44421 55873 44455
rect 55907 44452 55919 44455
rect 56318 44452 56324 44464
rect 55907 44424 56324 44452
rect 55907 44421 55919 44424
rect 55861 44415 55919 44421
rect 56318 44412 56324 44424
rect 56376 44452 56382 44464
rect 56689 44455 56747 44461
rect 56689 44452 56701 44455
rect 56376 44424 56701 44452
rect 56376 44412 56382 44424
rect 56689 44421 56701 44424
rect 56735 44421 56747 44455
rect 56689 44415 56747 44421
rect 54757 44387 54815 44393
rect 54757 44353 54769 44387
rect 54803 44384 54815 44387
rect 55398 44384 55404 44396
rect 54803 44356 55404 44384
rect 54803 44353 54815 44356
rect 54757 44347 54815 44353
rect 55398 44344 55404 44356
rect 55456 44384 55462 44396
rect 55677 44387 55735 44393
rect 55677 44384 55689 44387
rect 55456 44356 55689 44384
rect 55456 44344 55462 44356
rect 55677 44353 55689 44356
rect 55723 44353 55735 44387
rect 56502 44384 56508 44396
rect 56463 44356 56508 44384
rect 55677 44347 55735 44353
rect 56502 44344 56508 44356
rect 56560 44344 56566 44396
rect 56781 44387 56839 44393
rect 56781 44353 56793 44387
rect 56827 44384 56839 44387
rect 56962 44384 56968 44396
rect 56827 44356 56968 44384
rect 56827 44353 56839 44356
rect 56781 44347 56839 44353
rect 56962 44344 56968 44356
rect 57020 44344 57026 44396
rect 55306 44316 55312 44328
rect 54496 44288 55312 44316
rect 55306 44276 55312 44288
rect 55364 44316 55370 44328
rect 55585 44319 55643 44325
rect 55585 44316 55597 44319
rect 55364 44288 55597 44316
rect 55364 44276 55370 44288
rect 55585 44285 55597 44288
rect 55631 44285 55643 44319
rect 55585 44279 55643 44285
rect 55766 44276 55772 44328
rect 55824 44316 55830 44328
rect 56321 44319 56379 44325
rect 56321 44316 56333 44319
rect 55824 44288 56333 44316
rect 55824 44276 55830 44288
rect 56321 44285 56333 44288
rect 56367 44285 56379 44319
rect 56321 44279 56379 44285
rect 52144 44220 52960 44248
rect 52144 44208 52150 44220
rect 34885 44183 34943 44189
rect 34885 44180 34897 44183
rect 34572 44152 34897 44180
rect 34572 44140 34578 44152
rect 34885 44149 34897 44152
rect 34931 44149 34943 44183
rect 39666 44180 39672 44192
rect 39627 44152 39672 44180
rect 34885 44143 34943 44149
rect 39666 44140 39672 44152
rect 39724 44140 39730 44192
rect 42429 44183 42487 44189
rect 42429 44149 42441 44183
rect 42475 44180 42487 44183
rect 42794 44180 42800 44192
rect 42475 44152 42800 44180
rect 42475 44149 42487 44152
rect 42429 44143 42487 44149
rect 42794 44140 42800 44152
rect 42852 44140 42858 44192
rect 44913 44183 44971 44189
rect 44913 44149 44925 44183
rect 44959 44180 44971 44183
rect 46106 44180 46112 44192
rect 44959 44152 46112 44180
rect 44959 44149 44971 44152
rect 44913 44143 44971 44149
rect 46106 44140 46112 44152
rect 46164 44140 46170 44192
rect 46201 44183 46259 44189
rect 46201 44149 46213 44183
rect 46247 44180 46259 44183
rect 47670 44180 47676 44192
rect 46247 44152 47676 44180
rect 46247 44149 46259 44152
rect 46201 44143 46259 44149
rect 47670 44140 47676 44152
rect 47728 44140 47734 44192
rect 53098 44180 53104 44192
rect 53059 44152 53104 44180
rect 53098 44140 53104 44152
rect 53156 44140 53162 44192
rect 54478 44180 54484 44192
rect 54439 44152 54484 44180
rect 54478 44140 54484 44152
rect 54536 44140 54542 44192
rect 56594 44140 56600 44192
rect 56652 44180 56658 44192
rect 58069 44183 58127 44189
rect 58069 44180 58081 44183
rect 56652 44152 58081 44180
rect 56652 44140 56658 44152
rect 58069 44149 58081 44152
rect 58115 44149 58127 44183
rect 58069 44143 58127 44149
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 29454 43936 29460 43988
rect 29512 43976 29518 43988
rect 29549 43979 29607 43985
rect 29549 43976 29561 43979
rect 29512 43948 29561 43976
rect 29512 43936 29518 43948
rect 29549 43945 29561 43948
rect 29595 43945 29607 43979
rect 29549 43939 29607 43945
rect 35526 43936 35532 43988
rect 35584 43976 35590 43988
rect 35759 43979 35817 43985
rect 35759 43976 35771 43979
rect 35584 43948 35771 43976
rect 35584 43936 35590 43948
rect 35759 43945 35771 43948
rect 35805 43945 35817 43979
rect 35759 43939 35817 43945
rect 37550 43936 37556 43988
rect 37608 43976 37614 43988
rect 37737 43979 37795 43985
rect 37737 43976 37749 43979
rect 37608 43948 37749 43976
rect 37608 43936 37614 43948
rect 37737 43945 37749 43948
rect 37783 43945 37795 43979
rect 37737 43939 37795 43945
rect 38930 43936 38936 43988
rect 38988 43976 38994 43988
rect 39853 43979 39911 43985
rect 39853 43976 39865 43979
rect 38988 43948 39865 43976
rect 38988 43936 38994 43948
rect 39853 43945 39865 43948
rect 39899 43945 39911 43979
rect 39853 43939 39911 43945
rect 43073 43979 43131 43985
rect 43073 43945 43085 43979
rect 43119 43976 43131 43979
rect 43714 43976 43720 43988
rect 43119 43948 43720 43976
rect 43119 43945 43131 43948
rect 43073 43939 43131 43945
rect 43714 43936 43720 43948
rect 43772 43936 43778 43988
rect 44818 43936 44824 43988
rect 44876 43976 44882 43988
rect 44876 43948 45968 43976
rect 44876 43936 44882 43948
rect 32766 43868 32772 43920
rect 32824 43908 32830 43920
rect 39022 43908 39028 43920
rect 32824 43880 39028 43908
rect 32824 43868 32830 43880
rect 39022 43868 39028 43880
rect 39080 43868 39086 43920
rect 39114 43868 39120 43920
rect 39172 43908 39178 43920
rect 39209 43911 39267 43917
rect 39209 43908 39221 43911
rect 39172 43880 39221 43908
rect 39172 43868 39178 43880
rect 39209 43877 39221 43880
rect 39255 43877 39267 43911
rect 39209 43871 39267 43877
rect 39758 43868 39764 43920
rect 39816 43908 39822 43920
rect 39816 43880 42104 43908
rect 39816 43868 39822 43880
rect 27801 43843 27859 43849
rect 27801 43809 27813 43843
rect 27847 43840 27859 43843
rect 29086 43840 29092 43852
rect 27847 43812 29092 43840
rect 27847 43809 27859 43812
rect 27801 43803 27859 43809
rect 29086 43800 29092 43812
rect 29144 43800 29150 43852
rect 31018 43800 31024 43852
rect 31076 43840 31082 43852
rect 31113 43843 31171 43849
rect 31113 43840 31125 43843
rect 31076 43812 31125 43840
rect 31076 43800 31082 43812
rect 31113 43809 31125 43812
rect 31159 43809 31171 43843
rect 31113 43803 31171 43809
rect 38197 43843 38255 43849
rect 38197 43809 38209 43843
rect 38243 43840 38255 43843
rect 38841 43843 38899 43849
rect 38841 43840 38853 43843
rect 38243 43812 38853 43840
rect 38243 43809 38255 43812
rect 38197 43803 38255 43809
rect 38841 43809 38853 43812
rect 38887 43809 38899 43843
rect 40310 43840 40316 43852
rect 40271 43812 40316 43840
rect 38841 43803 38899 43809
rect 40310 43800 40316 43812
rect 40368 43800 40374 43852
rect 41966 43840 41972 43852
rect 41432 43812 41972 43840
rect 27985 43775 28043 43781
rect 27985 43741 27997 43775
rect 28031 43741 28043 43775
rect 27985 43735 28043 43741
rect 28169 43775 28227 43781
rect 28169 43741 28181 43775
rect 28215 43772 28227 43775
rect 29733 43775 29791 43781
rect 29733 43772 29745 43775
rect 28215 43744 29745 43772
rect 28215 43741 28227 43744
rect 28169 43735 28227 43741
rect 29733 43741 29745 43744
rect 29779 43741 29791 43775
rect 29733 43735 29791 43741
rect 31380 43775 31438 43781
rect 31380 43741 31392 43775
rect 31426 43772 31438 43775
rect 32122 43772 32128 43784
rect 31426 43744 32128 43772
rect 31426 43741 31438 43744
rect 31380 43735 31438 43741
rect 28000 43704 28028 43735
rect 32122 43732 32128 43744
rect 32180 43732 32186 43784
rect 35529 43775 35587 43781
rect 35529 43741 35541 43775
rect 35575 43772 35587 43775
rect 35894 43772 35900 43784
rect 35575 43744 35900 43772
rect 35575 43741 35587 43744
rect 35529 43735 35587 43741
rect 35894 43732 35900 43744
rect 35952 43732 35958 43784
rect 37921 43775 37979 43781
rect 37921 43741 37933 43775
rect 37967 43741 37979 43775
rect 37921 43735 37979 43741
rect 38013 43775 38071 43781
rect 38013 43741 38025 43775
rect 38059 43741 38071 43775
rect 38013 43735 38071 43741
rect 29086 43704 29092 43716
rect 28000 43676 29092 43704
rect 29086 43664 29092 43676
rect 29144 43664 29150 43716
rect 32398 43596 32404 43648
rect 32456 43636 32462 43648
rect 32493 43639 32551 43645
rect 32493 43636 32505 43639
rect 32456 43608 32505 43636
rect 32456 43596 32462 43608
rect 32493 43605 32505 43608
rect 32539 43605 32551 43639
rect 32493 43599 32551 43605
rect 34606 43596 34612 43648
rect 34664 43636 34670 43648
rect 35986 43636 35992 43648
rect 34664 43608 35992 43636
rect 34664 43596 34670 43608
rect 35986 43596 35992 43608
rect 36044 43596 36050 43648
rect 37936 43636 37964 43735
rect 38028 43704 38056 43735
rect 38102 43732 38108 43784
rect 38160 43772 38166 43784
rect 38746 43772 38752 43784
rect 38160 43744 38205 43772
rect 38707 43744 38752 43772
rect 38160 43732 38166 43744
rect 38746 43732 38752 43744
rect 38804 43732 38810 43784
rect 38930 43772 38936 43784
rect 38891 43744 38936 43772
rect 38930 43732 38936 43744
rect 38988 43732 38994 43784
rect 39025 43775 39083 43781
rect 39025 43741 39037 43775
rect 39071 43741 39083 43775
rect 39025 43735 39083 43741
rect 39301 43775 39359 43781
rect 39301 43741 39313 43775
rect 39347 43772 39359 43775
rect 39758 43772 39764 43784
rect 39347 43744 39764 43772
rect 39347 43741 39359 43744
rect 39301 43735 39359 43741
rect 38286 43704 38292 43716
rect 38028 43676 38292 43704
rect 38286 43664 38292 43676
rect 38344 43664 38350 43716
rect 38378 43664 38384 43716
rect 38436 43704 38442 43716
rect 39040 43704 39068 43735
rect 39758 43732 39764 43744
rect 39816 43732 39822 43784
rect 40034 43772 40040 43784
rect 39995 43744 40040 43772
rect 40034 43732 40040 43744
rect 40092 43732 40098 43784
rect 40129 43775 40187 43781
rect 40129 43741 40141 43775
rect 40175 43741 40187 43775
rect 40129 43735 40187 43741
rect 40405 43775 40463 43781
rect 40405 43741 40417 43775
rect 40451 43772 40463 43775
rect 40678 43772 40684 43784
rect 40451 43744 40684 43772
rect 40451 43741 40463 43744
rect 40405 43735 40463 43741
rect 40144 43704 40172 43735
rect 40678 43732 40684 43744
rect 40736 43732 40742 43784
rect 41138 43732 41144 43784
rect 41196 43772 41202 43784
rect 41432 43781 41460 43812
rect 41966 43800 41972 43812
rect 42024 43800 42030 43852
rect 42076 43840 42104 43880
rect 42150 43868 42156 43920
rect 42208 43908 42214 43920
rect 42521 43911 42579 43917
rect 42521 43908 42533 43911
rect 42208 43880 42533 43908
rect 42208 43868 42214 43880
rect 42521 43877 42533 43880
rect 42567 43877 42579 43911
rect 45554 43908 45560 43920
rect 42521 43871 42579 43877
rect 44008 43880 45560 43908
rect 44008 43840 44036 43880
rect 45554 43868 45560 43880
rect 45612 43868 45618 43920
rect 45940 43908 45968 43948
rect 46014 43936 46020 43988
rect 46072 43976 46078 43988
rect 46072 43948 50016 43976
rect 46072 43936 46078 43948
rect 45940 43880 46796 43908
rect 46768 43852 46796 43880
rect 46842 43868 46848 43920
rect 46900 43908 46906 43920
rect 47489 43911 47547 43917
rect 47489 43908 47501 43911
rect 46900 43880 47501 43908
rect 46900 43868 46906 43880
rect 47489 43877 47501 43880
rect 47535 43877 47547 43911
rect 47489 43871 47547 43877
rect 47581 43911 47639 43917
rect 47581 43877 47593 43911
rect 47627 43908 47639 43911
rect 48225 43911 48283 43917
rect 48225 43908 48237 43911
rect 47627 43880 48237 43908
rect 47627 43877 47639 43880
rect 47581 43871 47639 43877
rect 48225 43877 48237 43880
rect 48271 43908 48283 43911
rect 49326 43908 49332 43920
rect 48271 43880 49332 43908
rect 48271 43877 48283 43880
rect 48225 43871 48283 43877
rect 49326 43868 49332 43880
rect 49384 43868 49390 43920
rect 49988 43908 50016 43948
rect 50062 43936 50068 43988
rect 50120 43976 50126 43988
rect 50157 43979 50215 43985
rect 50157 43976 50169 43979
rect 50120 43948 50169 43976
rect 50120 43936 50126 43948
rect 50157 43945 50169 43948
rect 50203 43945 50215 43979
rect 52638 43976 52644 43988
rect 52599 43948 52644 43976
rect 50157 43939 50215 43945
rect 52638 43936 52644 43948
rect 52696 43936 52702 43988
rect 53834 43976 53840 43988
rect 53795 43948 53840 43976
rect 53834 43936 53840 43948
rect 53892 43936 53898 43988
rect 55122 43936 55128 43988
rect 55180 43976 55186 43988
rect 55493 43979 55551 43985
rect 55493 43976 55505 43979
rect 55180 43948 55505 43976
rect 55180 43936 55186 43948
rect 55493 43945 55505 43948
rect 55539 43945 55551 43979
rect 57146 43976 57152 43988
rect 55493 43939 55551 43945
rect 55600 43948 57152 43976
rect 55600 43908 55628 43948
rect 57146 43936 57152 43948
rect 57204 43936 57210 43988
rect 49988 43880 55628 43908
rect 55677 43911 55735 43917
rect 55677 43877 55689 43911
rect 55723 43877 55735 43911
rect 55677 43871 55735 43877
rect 44910 43840 44916 43852
rect 42076 43812 44036 43840
rect 44100 43812 44916 43840
rect 41325 43775 41383 43781
rect 41325 43772 41337 43775
rect 41196 43744 41337 43772
rect 41196 43732 41202 43744
rect 41325 43741 41337 43744
rect 41371 43741 41383 43775
rect 41325 43735 41383 43741
rect 41417 43775 41475 43781
rect 41417 43741 41429 43775
rect 41463 43741 41475 43775
rect 41601 43775 41659 43781
rect 41601 43772 41613 43775
rect 41417 43735 41475 43741
rect 41524 43744 41613 43772
rect 41046 43704 41052 43716
rect 38436 43676 41052 43704
rect 38436 43664 38442 43676
rect 41046 43664 41052 43676
rect 41104 43664 41110 43716
rect 40954 43636 40960 43648
rect 37936 43608 40960 43636
rect 40954 43596 40960 43608
rect 41012 43596 41018 43648
rect 41141 43639 41199 43645
rect 41141 43605 41153 43639
rect 41187 43636 41199 43639
rect 41322 43636 41328 43648
rect 41187 43608 41328 43636
rect 41187 43605 41199 43608
rect 41141 43599 41199 43605
rect 41322 43596 41328 43608
rect 41380 43596 41386 43648
rect 41524 43636 41552 43744
rect 41601 43741 41613 43744
rect 41647 43741 41659 43775
rect 41601 43735 41659 43741
rect 41703 43775 41761 43781
rect 41703 43741 41715 43775
rect 41749 43772 41761 43775
rect 42076 43772 42104 43812
rect 41749 43744 42104 43772
rect 41749 43741 41761 43744
rect 41703 43735 41761 43741
rect 42426 43732 42432 43784
rect 42484 43772 42490 43784
rect 44100 43781 44128 43812
rect 44910 43800 44916 43812
rect 44968 43800 44974 43852
rect 45186 43840 45192 43852
rect 45147 43812 45192 43840
rect 45186 43800 45192 43812
rect 45244 43800 45250 43852
rect 45646 43800 45652 43852
rect 45704 43800 45710 43852
rect 45738 43800 45744 43852
rect 45796 43840 45802 43852
rect 46661 43843 46719 43849
rect 46661 43840 46673 43843
rect 45796 43812 46673 43840
rect 45796 43800 45802 43812
rect 46661 43809 46673 43812
rect 46707 43809 46719 43843
rect 46661 43803 46719 43809
rect 46750 43800 46756 43852
rect 46808 43840 46814 43852
rect 49602 43840 49608 43852
rect 46808 43812 46901 43840
rect 47596 43812 49608 43840
rect 46808 43800 46814 43812
rect 44085 43775 44143 43781
rect 44085 43772 44097 43775
rect 42484 43744 44097 43772
rect 42484 43732 42490 43744
rect 44085 43741 44097 43744
rect 44131 43741 44143 43775
rect 44085 43735 44143 43741
rect 44174 43732 44180 43784
rect 44232 43772 44238 43784
rect 44361 43775 44419 43781
rect 44232 43744 44277 43772
rect 44232 43732 44238 43744
rect 44361 43741 44373 43775
rect 44407 43741 44419 43775
rect 44361 43735 44419 43741
rect 44453 43775 44511 43781
rect 44453 43741 44465 43775
rect 44499 43772 44511 43775
rect 45281 43775 45339 43781
rect 44499 43744 45140 43772
rect 44499 43741 44511 43744
rect 44453 43735 44511 43741
rect 42794 43704 42800 43716
rect 42755 43676 42800 43704
rect 42794 43664 42800 43676
rect 42852 43664 42858 43716
rect 42978 43664 42984 43716
rect 43036 43704 43042 43716
rect 43901 43707 43959 43713
rect 43901 43704 43913 43707
rect 43036 43676 43913 43704
rect 43036 43664 43042 43676
rect 43901 43673 43913 43676
rect 43947 43673 43959 43707
rect 44376 43704 44404 43735
rect 44910 43704 44916 43716
rect 44376 43676 44916 43704
rect 43901 43667 43959 43673
rect 44910 43664 44916 43676
rect 44968 43664 44974 43716
rect 41690 43636 41696 43648
rect 41524 43608 41696 43636
rect 41690 43596 41696 43608
rect 41748 43596 41754 43648
rect 42610 43596 42616 43648
rect 42668 43636 42674 43648
rect 42705 43639 42763 43645
rect 42705 43636 42717 43639
rect 42668 43608 42717 43636
rect 42668 43596 42674 43608
rect 42705 43605 42717 43608
rect 42751 43605 42763 43639
rect 42886 43636 42892 43648
rect 42847 43608 42892 43636
rect 42705 43599 42763 43605
rect 42886 43596 42892 43608
rect 42944 43596 42950 43648
rect 43990 43596 43996 43648
rect 44048 43636 44054 43648
rect 45005 43639 45063 43645
rect 45005 43636 45017 43639
rect 44048 43608 45017 43636
rect 44048 43596 44054 43608
rect 45005 43605 45017 43608
rect 45051 43605 45063 43639
rect 45112 43636 45140 43744
rect 45281 43741 45293 43775
rect 45327 43772 45339 43775
rect 45664 43772 45692 43800
rect 47596 43784 47624 43812
rect 49602 43800 49608 43812
rect 49660 43800 49666 43852
rect 50709 43843 50767 43849
rect 50709 43840 50721 43843
rect 50264 43812 50721 43840
rect 45327 43744 45692 43772
rect 46293 43775 46351 43781
rect 45327 43741 45339 43744
rect 45281 43735 45339 43741
rect 46293 43741 46305 43775
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 46385 43775 46443 43781
rect 46385 43741 46397 43775
rect 46431 43772 46443 43775
rect 46474 43772 46480 43784
rect 46431 43744 46480 43772
rect 46431 43741 46443 43744
rect 46385 43735 46443 43741
rect 45370 43664 45376 43716
rect 45428 43704 45434 43716
rect 45557 43707 45615 43713
rect 45557 43704 45569 43707
rect 45428 43676 45569 43704
rect 45428 43664 45434 43676
rect 45557 43673 45569 43676
rect 45603 43673 45615 43707
rect 45557 43667 45615 43673
rect 45646 43664 45652 43716
rect 45704 43704 45710 43716
rect 46308 43704 46336 43735
rect 46474 43732 46480 43744
rect 46532 43732 46538 43784
rect 47397 43775 47455 43781
rect 47397 43741 47409 43775
rect 47443 43772 47455 43775
rect 47578 43772 47584 43784
rect 47443 43744 47584 43772
rect 47443 43741 47455 43744
rect 47397 43735 47455 43741
rect 47578 43732 47584 43744
rect 47636 43732 47642 43784
rect 47673 43775 47731 43781
rect 47673 43741 47685 43775
rect 47719 43741 47731 43775
rect 47673 43735 47731 43741
rect 47688 43704 47716 43735
rect 48130 43732 48136 43784
rect 48188 43772 48194 43784
rect 48225 43775 48283 43781
rect 48225 43772 48237 43775
rect 48188 43744 48237 43772
rect 48188 43732 48194 43744
rect 48225 43741 48237 43744
rect 48271 43741 48283 43775
rect 48225 43735 48283 43741
rect 48409 43775 48467 43781
rect 48409 43741 48421 43775
rect 48455 43772 48467 43775
rect 48590 43772 48596 43784
rect 48455 43744 48596 43772
rect 48455 43741 48467 43744
rect 48409 43735 48467 43741
rect 48590 43732 48596 43744
rect 48648 43732 48654 43784
rect 50062 43732 50068 43784
rect 50120 43772 50126 43784
rect 50264 43772 50292 43812
rect 50709 43809 50721 43812
rect 50755 43840 50767 43843
rect 50982 43840 50988 43852
rect 50755 43812 50988 43840
rect 50755 43809 50767 43812
rect 50709 43803 50767 43809
rect 50982 43800 50988 43812
rect 51040 43800 51046 43852
rect 52365 43843 52423 43849
rect 52365 43809 52377 43843
rect 52411 43809 52423 43843
rect 55692 43840 55720 43871
rect 52365 43803 52423 43809
rect 54404 43812 55720 43840
rect 56321 43843 56379 43849
rect 50120 43744 50292 43772
rect 50338 43775 50396 43781
rect 50120 43732 50126 43744
rect 50338 43741 50350 43775
rect 50384 43772 50396 43775
rect 50614 43772 50620 43784
rect 50384 43744 50620 43772
rect 50384 43741 50396 43744
rect 50338 43735 50396 43741
rect 50614 43732 50620 43744
rect 50672 43732 50678 43784
rect 50798 43732 50804 43784
rect 50856 43772 50862 43784
rect 52270 43772 52276 43784
rect 50856 43744 50901 43772
rect 52231 43744 52276 43772
rect 50856 43732 50862 43744
rect 52270 43732 52276 43744
rect 52328 43732 52334 43784
rect 52380 43772 52408 43803
rect 52914 43772 52920 43784
rect 52380 43744 52920 43772
rect 52914 43732 52920 43744
rect 52972 43732 52978 43784
rect 53745 43775 53803 43781
rect 53745 43741 53757 43775
rect 53791 43772 53803 43775
rect 53834 43772 53840 43784
rect 53791 43744 53840 43772
rect 53791 43741 53803 43744
rect 53745 43735 53803 43741
rect 53834 43732 53840 43744
rect 53892 43732 53898 43784
rect 53929 43775 53987 43781
rect 53929 43741 53941 43775
rect 53975 43772 53987 43775
rect 54294 43772 54300 43784
rect 53975 43744 54300 43772
rect 53975 43741 53987 43744
rect 53929 43735 53987 43741
rect 54294 43732 54300 43744
rect 54352 43732 54358 43784
rect 54404 43781 54432 43812
rect 56321 43809 56333 43843
rect 56367 43840 56379 43843
rect 56594 43840 56600 43852
rect 56367 43812 56600 43840
rect 56367 43809 56379 43812
rect 56321 43803 56379 43809
rect 56594 43800 56600 43812
rect 56652 43800 56658 43852
rect 57882 43840 57888 43852
rect 57843 43812 57888 43840
rect 57882 43800 57888 43812
rect 57940 43800 57946 43852
rect 54389 43775 54447 43781
rect 54389 43741 54401 43775
rect 54435 43741 54447 43775
rect 54389 43735 54447 43741
rect 54478 43732 54484 43784
rect 54536 43772 54542 43784
rect 54573 43775 54631 43781
rect 54573 43772 54585 43775
rect 54536 43744 54585 43772
rect 54536 43732 54542 43744
rect 54573 43741 54585 43744
rect 54619 43741 54631 43775
rect 54573 43735 54631 43741
rect 55306 43704 55312 43716
rect 45704 43676 46336 43704
rect 46860 43676 47716 43704
rect 55267 43676 55312 43704
rect 45704 43664 45710 43676
rect 46109 43639 46167 43645
rect 46109 43636 46121 43639
rect 45112 43608 46121 43636
rect 45005 43599 45063 43605
rect 46109 43605 46121 43608
rect 46155 43605 46167 43639
rect 46109 43599 46167 43605
rect 46198 43596 46204 43648
rect 46256 43636 46262 43648
rect 46860 43636 46888 43676
rect 55306 43664 55312 43676
rect 55364 43664 55370 43716
rect 55950 43664 55956 43716
rect 56008 43704 56014 43716
rect 56505 43707 56563 43713
rect 56505 43704 56517 43707
rect 56008 43676 56517 43704
rect 56008 43664 56014 43676
rect 56505 43673 56517 43676
rect 56551 43673 56563 43707
rect 56505 43667 56563 43673
rect 46256 43608 46888 43636
rect 47213 43639 47271 43645
rect 46256 43596 46262 43608
rect 47213 43605 47225 43639
rect 47259 43636 47271 43639
rect 47854 43636 47860 43648
rect 47259 43608 47860 43636
rect 47259 43605 47271 43608
rect 47213 43599 47271 43605
rect 47854 43596 47860 43608
rect 47912 43596 47918 43648
rect 50341 43639 50399 43645
rect 50341 43605 50353 43639
rect 50387 43636 50399 43639
rect 50614 43636 50620 43648
rect 50387 43608 50620 43636
rect 50387 43605 50399 43608
rect 50341 43599 50399 43605
rect 50614 43596 50620 43608
rect 50672 43596 50678 43648
rect 54754 43636 54760 43648
rect 54715 43608 54760 43636
rect 54754 43596 54760 43608
rect 54812 43596 54818 43648
rect 55398 43596 55404 43648
rect 55456 43636 55462 43648
rect 55509 43639 55567 43645
rect 55509 43636 55521 43639
rect 55456 43608 55521 43636
rect 55456 43596 55462 43608
rect 55509 43605 55521 43608
rect 55555 43605 55567 43639
rect 55509 43599 55567 43605
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 25501 43435 25559 43441
rect 25501 43401 25513 43435
rect 25547 43401 25559 43435
rect 41322 43432 41328 43444
rect 25501 43395 25559 43401
rect 35084 43404 41184 43432
rect 41283 43404 41328 43432
rect 24210 43324 24216 43376
rect 24268 43364 24274 43376
rect 25317 43367 25375 43373
rect 25317 43364 25329 43367
rect 24268 43336 25329 43364
rect 24268 43324 24274 43336
rect 25317 43333 25329 43336
rect 25363 43333 25375 43367
rect 25516 43364 25544 43395
rect 26234 43364 26240 43376
rect 25516 43336 26240 43364
rect 25317 43327 25375 43333
rect 26234 43324 26240 43336
rect 26292 43364 26298 43376
rect 26292 43336 26464 43364
rect 26292 43324 26298 43336
rect 22281 43299 22339 43305
rect 22281 43265 22293 43299
rect 22327 43265 22339 43299
rect 22281 43259 22339 43265
rect 23109 43299 23167 43305
rect 23109 43265 23121 43299
rect 23155 43296 23167 43299
rect 23290 43296 23296 43308
rect 23155 43268 23296 43296
rect 23155 43265 23167 43268
rect 23109 43259 23167 43265
rect 22296 43228 22324 43259
rect 23290 43256 23296 43268
rect 23348 43296 23354 43308
rect 24121 43299 24179 43305
rect 23348 43268 23704 43296
rect 23348 43256 23354 43268
rect 23676 43228 23704 43268
rect 24121 43265 24133 43299
rect 24167 43296 24179 43299
rect 25222 43296 25228 43308
rect 24167 43268 25228 43296
rect 24167 43265 24179 43268
rect 24121 43259 24179 43265
rect 25222 43256 25228 43268
rect 25280 43256 25286 43308
rect 26050 43256 26056 43308
rect 26108 43296 26114 43308
rect 26145 43299 26203 43305
rect 26145 43296 26157 43299
rect 26108 43268 26157 43296
rect 26108 43256 26114 43268
rect 26145 43265 26157 43268
rect 26191 43265 26203 43299
rect 26326 43296 26332 43308
rect 26287 43268 26332 43296
rect 26145 43259 26203 43265
rect 26326 43256 26332 43268
rect 26384 43256 26390 43308
rect 26436 43305 26464 43336
rect 26421 43299 26479 43305
rect 26421 43265 26433 43299
rect 26467 43265 26479 43299
rect 26421 43259 26479 43265
rect 34606 43256 34612 43308
rect 34664 43296 34670 43308
rect 35084 43305 35112 43404
rect 38657 43367 38715 43373
rect 38657 43364 38669 43367
rect 36188 43336 38669 43364
rect 34793 43299 34851 43305
rect 34793 43296 34805 43299
rect 34664 43268 34805 43296
rect 34664 43256 34670 43268
rect 34793 43265 34805 43268
rect 34839 43265 34851 43299
rect 34793 43259 34851 43265
rect 34977 43299 35035 43305
rect 34977 43265 34989 43299
rect 35023 43265 35035 43299
rect 34977 43259 35035 43265
rect 35069 43299 35127 43305
rect 35069 43265 35081 43299
rect 35115 43265 35127 43299
rect 35069 43259 35127 43265
rect 35345 43299 35403 43305
rect 35345 43265 35357 43299
rect 35391 43296 35403 43299
rect 35526 43296 35532 43308
rect 35391 43268 35532 43296
rect 35391 43265 35403 43268
rect 35345 43259 35403 43265
rect 24213 43231 24271 43237
rect 24213 43228 24225 43231
rect 22296 43200 23520 43228
rect 23676 43200 24225 43228
rect 23492 43172 23520 43200
rect 24213 43197 24225 43200
rect 24259 43197 24271 43231
rect 24213 43191 24271 43197
rect 24305 43231 24363 43237
rect 24305 43197 24317 43231
rect 24351 43197 24363 43231
rect 24305 43191 24363 43197
rect 23474 43120 23480 43172
rect 23532 43160 23538 43172
rect 24320 43160 24348 43191
rect 24394 43188 24400 43240
rect 24452 43228 24458 43240
rect 24452 43200 24497 43228
rect 24452 43188 24458 43200
rect 23532 43132 24348 43160
rect 23532 43120 23538 43132
rect 24486 43120 24492 43172
rect 24544 43160 24550 43172
rect 24949 43163 25007 43169
rect 24949 43160 24961 43163
rect 24544 43132 24961 43160
rect 24544 43120 24550 43132
rect 24949 43129 24961 43132
rect 24995 43129 25007 43163
rect 34992 43160 35020 43259
rect 35526 43256 35532 43268
rect 35584 43296 35590 43308
rect 35584 43268 35940 43296
rect 35584 43256 35590 43268
rect 35161 43231 35219 43237
rect 35161 43197 35173 43231
rect 35207 43228 35219 43231
rect 35618 43228 35624 43240
rect 35207 43200 35624 43228
rect 35207 43197 35219 43200
rect 35161 43191 35219 43197
rect 35618 43188 35624 43200
rect 35676 43188 35682 43240
rect 35434 43160 35440 43172
rect 34992 43132 35440 43160
rect 24949 43123 25007 43129
rect 35434 43120 35440 43132
rect 35492 43120 35498 43172
rect 35912 43160 35940 43268
rect 35986 43256 35992 43308
rect 36044 43296 36050 43308
rect 36188 43305 36216 43336
rect 38657 43333 38669 43336
rect 38703 43333 38715 43367
rect 41156 43364 41184 43404
rect 41322 43392 41328 43404
rect 41380 43392 41386 43444
rect 42610 43392 42616 43444
rect 42668 43432 42674 43444
rect 42794 43432 42800 43444
rect 42668 43404 42800 43432
rect 42668 43392 42674 43404
rect 42794 43392 42800 43404
rect 42852 43392 42858 43444
rect 42886 43392 42892 43444
rect 42944 43432 42950 43444
rect 43165 43435 43223 43441
rect 43165 43432 43177 43435
rect 42944 43404 43177 43432
rect 42944 43392 42950 43404
rect 43165 43401 43177 43404
rect 43211 43401 43223 43435
rect 43165 43395 43223 43401
rect 43717 43435 43775 43441
rect 43717 43401 43729 43435
rect 43763 43401 43775 43435
rect 43717 43395 43775 43401
rect 43732 43364 43760 43395
rect 44634 43392 44640 43444
rect 44692 43432 44698 43444
rect 44729 43435 44787 43441
rect 44729 43432 44741 43435
rect 44692 43404 44741 43432
rect 44692 43392 44698 43404
rect 44729 43401 44741 43404
rect 44775 43432 44787 43435
rect 45554 43432 45560 43444
rect 44775 43404 45560 43432
rect 44775 43401 44787 43404
rect 44729 43395 44787 43401
rect 45554 43392 45560 43404
rect 45612 43392 45618 43444
rect 46017 43435 46075 43441
rect 46017 43401 46029 43435
rect 46063 43432 46075 43435
rect 46198 43432 46204 43444
rect 46063 43404 46204 43432
rect 46063 43401 46075 43404
rect 46017 43395 46075 43401
rect 46198 43392 46204 43404
rect 46256 43392 46262 43444
rect 46474 43432 46480 43444
rect 46435 43404 46480 43432
rect 46474 43392 46480 43404
rect 46532 43392 46538 43444
rect 46934 43392 46940 43444
rect 46992 43432 46998 43444
rect 47210 43432 47216 43444
rect 46992 43404 47216 43432
rect 46992 43392 46998 43404
rect 47210 43392 47216 43404
rect 47268 43392 47274 43444
rect 50706 43432 50712 43444
rect 50667 43404 50712 43432
rect 50706 43392 50712 43404
rect 50764 43392 50770 43444
rect 50798 43392 50804 43444
rect 50856 43432 50862 43444
rect 51629 43435 51687 43441
rect 51629 43432 51641 43435
rect 50856 43404 51641 43432
rect 50856 43392 50862 43404
rect 51629 43401 51641 43404
rect 51675 43401 51687 43435
rect 54294 43432 54300 43444
rect 54255 43404 54300 43432
rect 51629 43395 51687 43401
rect 54294 43392 54300 43404
rect 54352 43392 54358 43444
rect 55122 43432 55128 43444
rect 55083 43404 55128 43432
rect 55122 43392 55128 43404
rect 55180 43392 55186 43444
rect 55493 43435 55551 43441
rect 55493 43401 55505 43435
rect 55539 43432 55551 43435
rect 55582 43432 55588 43444
rect 55539 43404 55588 43432
rect 55539 43401 55551 43404
rect 55493 43395 55551 43401
rect 55582 43392 55588 43404
rect 55640 43392 55646 43444
rect 57146 43432 57152 43444
rect 57107 43404 57152 43432
rect 57146 43392 57152 43404
rect 57204 43392 57210 43444
rect 41156 43336 43760 43364
rect 43809 43367 43867 43373
rect 38657 43327 38715 43333
rect 43809 43333 43821 43367
rect 43855 43364 43867 43367
rect 44361 43367 44419 43373
rect 44361 43364 44373 43367
rect 43855 43336 44373 43364
rect 43855 43333 43867 43336
rect 43809 43327 43867 43333
rect 44361 43333 44373 43336
rect 44407 43333 44419 43367
rect 44361 43327 44419 43333
rect 44468 43336 44864 43364
rect 36173 43299 36231 43305
rect 36044 43268 36089 43296
rect 36044 43256 36050 43268
rect 36173 43265 36185 43299
rect 36219 43265 36231 43299
rect 36173 43259 36231 43265
rect 36262 43256 36268 43308
rect 36320 43296 36326 43308
rect 36541 43299 36599 43305
rect 36320 43268 36365 43296
rect 36320 43256 36326 43268
rect 36541 43265 36553 43299
rect 36587 43265 36599 43299
rect 38378 43296 38384 43308
rect 38339 43268 38384 43296
rect 36541 43259 36599 43265
rect 36078 43188 36084 43240
rect 36136 43228 36142 43240
rect 36357 43231 36415 43237
rect 36357 43228 36369 43231
rect 36136 43200 36369 43228
rect 36136 43188 36142 43200
rect 36357 43197 36369 43200
rect 36403 43197 36415 43231
rect 36357 43191 36415 43197
rect 36556 43160 36584 43259
rect 38378 43256 38384 43268
rect 38436 43256 38442 43308
rect 41230 43296 41236 43308
rect 41191 43268 41236 43296
rect 41230 43256 41236 43268
rect 41288 43256 41294 43308
rect 41417 43299 41475 43305
rect 41417 43265 41429 43299
rect 41463 43265 41475 43299
rect 41417 43259 41475 43265
rect 38657 43231 38715 43237
rect 38657 43197 38669 43231
rect 38703 43228 38715 43231
rect 40957 43231 41015 43237
rect 40957 43228 40969 43231
rect 38703 43200 40969 43228
rect 38703 43197 38715 43200
rect 38657 43191 38715 43197
rect 40957 43197 40969 43200
rect 41003 43197 41015 43231
rect 40957 43191 41015 43197
rect 35912 43132 36584 43160
rect 22554 43092 22560 43104
rect 22515 43064 22560 43092
rect 22554 43052 22560 43064
rect 22612 43052 22618 43104
rect 23293 43095 23351 43101
rect 23293 43061 23305 43095
rect 23339 43092 23351 43095
rect 23382 43092 23388 43104
rect 23339 43064 23388 43092
rect 23339 43061 23351 43064
rect 23293 43055 23351 43061
rect 23382 43052 23388 43064
rect 23440 43052 23446 43104
rect 23937 43095 23995 43101
rect 23937 43061 23949 43095
rect 23983 43092 23995 43095
rect 24670 43092 24676 43104
rect 23983 43064 24676 43092
rect 23983 43061 23995 43064
rect 23937 43055 23995 43061
rect 24670 43052 24676 43064
rect 24728 43092 24734 43104
rect 25317 43095 25375 43101
rect 25317 43092 25329 43095
rect 24728 43064 25329 43092
rect 24728 43052 24734 43064
rect 25317 43061 25329 43064
rect 25363 43061 25375 43095
rect 25958 43092 25964 43104
rect 25919 43064 25964 43092
rect 25317 43055 25375 43061
rect 25958 43052 25964 43064
rect 26016 43052 26022 43104
rect 35526 43092 35532 43104
rect 35487 43064 35532 43092
rect 35526 43052 35532 43064
rect 35584 43052 35590 43104
rect 36722 43092 36728 43104
rect 36683 43064 36728 43092
rect 36722 43052 36728 43064
rect 36780 43052 36786 43104
rect 37734 43052 37740 43104
rect 37792 43092 37798 43104
rect 38473 43095 38531 43101
rect 38473 43092 38485 43095
rect 37792 43064 38485 43092
rect 37792 43052 37798 43064
rect 38473 43061 38485 43064
rect 38519 43061 38531 43095
rect 38473 43055 38531 43061
rect 40954 43052 40960 43104
rect 41012 43092 41018 43104
rect 41432 43092 41460 43259
rect 41782 43256 41788 43308
rect 41840 43296 41846 43308
rect 42429 43299 42487 43305
rect 42429 43296 42441 43299
rect 41840 43268 42441 43296
rect 41840 43256 41846 43268
rect 42429 43265 42441 43268
rect 42475 43265 42487 43299
rect 42429 43259 42487 43265
rect 42518 43256 42524 43308
rect 42576 43296 42582 43308
rect 42613 43299 42671 43305
rect 42613 43296 42625 43299
rect 42576 43268 42625 43296
rect 42576 43256 42582 43268
rect 42613 43265 42625 43268
rect 42659 43265 42671 43299
rect 42613 43259 42671 43265
rect 42705 43299 42763 43305
rect 42705 43265 42717 43299
rect 42751 43296 42763 43299
rect 42886 43296 42892 43308
rect 42751 43268 42892 43296
rect 42751 43265 42763 43268
rect 42705 43259 42763 43265
rect 42886 43256 42892 43268
rect 42944 43256 42950 43308
rect 42981 43299 43039 43305
rect 42981 43265 42993 43299
rect 43027 43296 43039 43299
rect 43162 43296 43168 43308
rect 43027 43268 43168 43296
rect 43027 43265 43039 43268
rect 42981 43259 43039 43265
rect 43162 43256 43168 43268
rect 43220 43256 43226 43308
rect 43625 43299 43683 43305
rect 43625 43265 43637 43299
rect 43671 43265 43683 43299
rect 43625 43259 43683 43265
rect 43901 43299 43959 43305
rect 43901 43265 43913 43299
rect 43947 43296 43959 43299
rect 43990 43296 43996 43308
rect 43947 43268 43996 43296
rect 43947 43265 43959 43268
rect 43901 43259 43959 43265
rect 41693 43231 41751 43237
rect 41693 43197 41705 43231
rect 41739 43228 41751 43231
rect 42150 43228 42156 43240
rect 41739 43200 42156 43228
rect 41739 43197 41751 43200
rect 41693 43191 41751 43197
rect 42150 43188 42156 43200
rect 42208 43188 42214 43240
rect 42242 43188 42248 43240
rect 42300 43228 42306 43240
rect 42797 43231 42855 43237
rect 42797 43228 42809 43231
rect 42300 43200 42809 43228
rect 42300 43188 42306 43200
rect 42797 43197 42809 43200
rect 42843 43197 42855 43231
rect 43640 43228 43668 43259
rect 43990 43256 43996 43268
rect 44048 43256 44054 43308
rect 44082 43256 44088 43308
rect 44140 43296 44146 43308
rect 44468 43296 44496 43336
rect 44836 43305 44864 43336
rect 44910 43324 44916 43376
rect 44968 43364 44974 43376
rect 47857 43367 47915 43373
rect 47857 43364 47869 43367
rect 44968 43336 47869 43364
rect 44968 43324 44974 43336
rect 47857 43333 47869 43336
rect 47903 43333 47915 43367
rect 54312 43364 54340 43392
rect 54312 43336 55628 43364
rect 47857 43327 47915 43333
rect 44140 43268 44496 43296
rect 44545 43299 44603 43305
rect 44140 43256 44146 43268
rect 44545 43265 44557 43299
rect 44591 43265 44603 43299
rect 44545 43259 44603 43265
rect 44821 43299 44879 43305
rect 44821 43265 44833 43299
rect 44867 43265 44879 43299
rect 44821 43259 44879 43265
rect 44450 43228 44456 43240
rect 43640 43200 44456 43228
rect 42797 43191 42855 43197
rect 42812 43160 42840 43191
rect 44450 43188 44456 43200
rect 44508 43188 44514 43240
rect 43070 43160 43076 43172
rect 42812 43132 43076 43160
rect 43070 43120 43076 43132
rect 43128 43120 43134 43172
rect 41012 43064 41460 43092
rect 41601 43095 41659 43101
rect 41012 43052 41018 43064
rect 41601 43061 41613 43095
rect 41647 43092 41659 43095
rect 44266 43092 44272 43104
rect 41647 43064 44272 43092
rect 41647 43061 41659 43064
rect 41601 43055 41659 43061
rect 44266 43052 44272 43064
rect 44324 43052 44330 43104
rect 44560 43092 44588 43259
rect 44836 43160 44864 43259
rect 45002 43256 45008 43308
rect 45060 43296 45066 43308
rect 45281 43299 45339 43305
rect 45281 43296 45293 43299
rect 45060 43268 45293 43296
rect 45060 43256 45066 43268
rect 45281 43265 45293 43268
rect 45327 43265 45339 43299
rect 45462 43296 45468 43308
rect 45423 43268 45468 43296
rect 45281 43259 45339 43265
rect 45462 43256 45468 43268
rect 45520 43256 45526 43308
rect 45554 43256 45560 43308
rect 45612 43296 45618 43308
rect 45830 43296 45836 43308
rect 45612 43268 45657 43296
rect 45791 43268 45836 43296
rect 45612 43256 45618 43268
rect 45830 43256 45836 43268
rect 45888 43256 45894 43308
rect 46566 43256 46572 43308
rect 46624 43296 46630 43308
rect 46661 43299 46719 43305
rect 46661 43296 46673 43299
rect 46624 43268 46673 43296
rect 46624 43256 46630 43268
rect 46661 43265 46673 43268
rect 46707 43265 46719 43299
rect 46661 43259 46719 43265
rect 47486 43256 47492 43308
rect 47544 43296 47550 43308
rect 47581 43299 47639 43305
rect 47581 43296 47593 43299
rect 47544 43268 47593 43296
rect 47544 43256 47550 43268
rect 47581 43265 47593 43268
rect 47627 43265 47639 43299
rect 47581 43259 47639 43265
rect 47670 43256 47676 43308
rect 47728 43296 47734 43308
rect 49053 43299 49111 43305
rect 47728 43268 47773 43296
rect 47728 43256 47734 43268
rect 49053 43265 49065 43299
rect 49099 43296 49111 43299
rect 49970 43296 49976 43308
rect 49099 43268 49976 43296
rect 49099 43265 49111 43268
rect 49053 43259 49111 43265
rect 49970 43256 49976 43268
rect 50028 43256 50034 43308
rect 50826 43299 50884 43305
rect 50826 43265 50838 43299
rect 50872 43296 50884 43299
rect 51442 43296 51448 43308
rect 50872 43268 51448 43296
rect 50872 43265 50884 43268
rect 50826 43259 50884 43265
rect 51442 43256 51448 43268
rect 51500 43256 51506 43308
rect 52270 43256 52276 43308
rect 52328 43296 52334 43308
rect 52733 43299 52791 43305
rect 52733 43296 52745 43299
rect 52328 43268 52745 43296
rect 52328 43256 52334 43268
rect 52733 43265 52745 43268
rect 52779 43265 52791 43299
rect 52914 43296 52920 43308
rect 52875 43268 52920 43296
rect 52733 43259 52791 43265
rect 52914 43256 52920 43268
rect 52972 43256 52978 43308
rect 53098 43256 53104 43308
rect 53156 43296 53162 43308
rect 53193 43299 53251 43305
rect 53193 43296 53205 43299
rect 53156 43268 53205 43296
rect 53156 43256 53162 43268
rect 53193 43265 53205 43268
rect 53239 43265 53251 43299
rect 53466 43296 53472 43308
rect 53427 43268 53472 43296
rect 53193 43259 53251 43265
rect 53466 43256 53472 43268
rect 53524 43256 53530 43308
rect 54018 43256 54024 43308
rect 54076 43296 54082 43308
rect 54205 43299 54263 43305
rect 54205 43296 54217 43299
rect 54076 43268 54217 43296
rect 54076 43256 54082 43268
rect 54205 43265 54217 43268
rect 54251 43265 54263 43299
rect 54386 43296 54392 43308
rect 54347 43268 54392 43296
rect 54205 43259 54263 43265
rect 54386 43256 54392 43268
rect 54444 43256 54450 43308
rect 55306 43296 55312 43308
rect 55267 43268 55312 43296
rect 55306 43256 55312 43268
rect 55364 43256 55370 43308
rect 55490 43256 55496 43308
rect 55548 43296 55554 43308
rect 55600 43305 55628 43336
rect 55585 43299 55643 43305
rect 55585 43296 55597 43299
rect 55548 43268 55597 43296
rect 55548 43256 55554 43268
rect 55585 43265 55597 43268
rect 55631 43265 55643 43299
rect 56318 43296 56324 43308
rect 56279 43268 56324 43296
rect 55585 43259 55643 43265
rect 56318 43256 56324 43268
rect 56376 43256 56382 43308
rect 57698 43256 57704 43308
rect 57756 43296 57762 43308
rect 57885 43299 57943 43305
rect 57885 43296 57897 43299
rect 57756 43268 57897 43296
rect 57756 43256 57762 43268
rect 57885 43265 57897 43268
rect 57931 43265 57943 43299
rect 57885 43259 57943 43265
rect 45186 43188 45192 43240
rect 45244 43228 45250 43240
rect 45649 43231 45707 43237
rect 45649 43228 45661 43231
rect 45244 43200 45661 43228
rect 45244 43188 45250 43200
rect 45649 43197 45661 43200
rect 45695 43197 45707 43231
rect 45649 43191 45707 43197
rect 46382 43188 46388 43240
rect 46440 43228 46446 43240
rect 46845 43231 46903 43237
rect 46845 43228 46857 43231
rect 46440 43200 46857 43228
rect 46440 43188 46446 43200
rect 46845 43197 46857 43200
rect 46891 43197 46903 43231
rect 46845 43191 46903 43197
rect 46937 43231 46995 43237
rect 46937 43197 46949 43231
rect 46983 43228 46995 43231
rect 47210 43228 47216 43240
rect 46983 43200 47216 43228
rect 46983 43197 46995 43200
rect 46937 43191 46995 43197
rect 47210 43188 47216 43200
rect 47268 43188 47274 43240
rect 47854 43228 47860 43240
rect 47815 43200 47860 43228
rect 47854 43188 47860 43200
rect 47912 43188 47918 43240
rect 49329 43231 49387 43237
rect 49329 43228 49341 43231
rect 48286 43200 49341 43228
rect 44836 43132 46980 43160
rect 46952 43104 46980 43132
rect 47302 43120 47308 43172
rect 47360 43160 47366 43172
rect 48130 43160 48136 43172
rect 47360 43132 48136 43160
rect 47360 43120 47366 43132
rect 48130 43120 48136 43132
rect 48188 43160 48194 43172
rect 48286 43160 48314 43200
rect 49329 43197 49341 43200
rect 49375 43197 49387 43231
rect 49329 43191 49387 43197
rect 50062 43188 50068 43240
rect 50120 43228 50126 43240
rect 50341 43231 50399 43237
rect 50341 43228 50353 43231
rect 50120 43200 50353 43228
rect 50120 43188 50126 43200
rect 50341 43197 50353 43200
rect 50387 43197 50399 43231
rect 50614 43228 50620 43240
rect 50575 43200 50620 43228
rect 50341 43191 50399 43197
rect 50614 43188 50620 43200
rect 50672 43188 50678 43240
rect 56505 43231 56563 43237
rect 56505 43197 56517 43231
rect 56551 43228 56563 43231
rect 56962 43228 56968 43240
rect 56551 43200 56968 43228
rect 56551 43197 56563 43200
rect 56505 43191 56563 43197
rect 56962 43188 56968 43200
rect 57020 43188 57026 43240
rect 48188 43132 48314 43160
rect 48188 43120 48194 43132
rect 50890 43120 50896 43172
rect 50948 43160 50954 43172
rect 50985 43163 51043 43169
rect 50985 43160 50997 43163
rect 50948 43132 50997 43160
rect 50948 43120 50954 43132
rect 50985 43129 50997 43132
rect 51031 43129 51043 43163
rect 50985 43123 51043 43129
rect 53101 43163 53159 43169
rect 53101 43129 53113 43163
rect 53147 43160 53159 43163
rect 54110 43160 54116 43172
rect 53147 43132 54116 43160
rect 53147 43129 53159 43132
rect 53101 43123 53159 43129
rect 54110 43120 54116 43132
rect 54168 43120 54174 43172
rect 45922 43092 45928 43104
rect 44560 43064 45928 43092
rect 45922 43052 45928 43064
rect 45980 43092 45986 43104
rect 46474 43092 46480 43104
rect 45980 43064 46480 43092
rect 45980 43052 45986 43064
rect 46474 43052 46480 43064
rect 46532 43052 46538 43104
rect 46934 43052 46940 43104
rect 46992 43052 46998 43104
rect 56870 43052 56876 43104
rect 56928 43092 56934 43104
rect 57977 43095 58035 43101
rect 57977 43092 57989 43095
rect 56928 43064 57989 43092
rect 56928 43052 56934 43064
rect 57977 43061 57989 43064
rect 58023 43061 58035 43095
rect 57977 43055 58035 43061
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 21450 42848 21456 42900
rect 21508 42888 21514 42900
rect 23382 42888 23388 42900
rect 21508 42860 23388 42888
rect 21508 42848 21514 42860
rect 23382 42848 23388 42860
rect 23440 42888 23446 42900
rect 33410 42888 33416 42900
rect 23440 42860 33416 42888
rect 23440 42848 23446 42860
rect 33410 42848 33416 42860
rect 33468 42848 33474 42900
rect 37734 42888 37740 42900
rect 37695 42860 37740 42888
rect 37734 42848 37740 42860
rect 37792 42848 37798 42900
rect 38749 42891 38807 42897
rect 38749 42857 38761 42891
rect 38795 42888 38807 42891
rect 40034 42888 40040 42900
rect 38795 42860 40040 42888
rect 38795 42857 38807 42860
rect 38749 42851 38807 42857
rect 40034 42848 40040 42860
rect 40092 42848 40098 42900
rect 41230 42848 41236 42900
rect 41288 42888 41294 42900
rect 41325 42891 41383 42897
rect 41325 42888 41337 42891
rect 41288 42860 41337 42888
rect 41288 42848 41294 42860
rect 41325 42857 41337 42860
rect 41371 42857 41383 42891
rect 42242 42888 42248 42900
rect 41325 42851 41383 42857
rect 41984 42860 42248 42888
rect 22557 42823 22615 42829
rect 22557 42789 22569 42823
rect 22603 42820 22615 42823
rect 22738 42820 22744 42832
rect 22603 42792 22744 42820
rect 22603 42789 22615 42792
rect 22557 42783 22615 42789
rect 22738 42780 22744 42792
rect 22796 42820 22802 42832
rect 23290 42820 23296 42832
rect 22796 42792 23296 42820
rect 22796 42780 22802 42792
rect 23290 42780 23296 42792
rect 23348 42820 23354 42832
rect 23569 42823 23627 42829
rect 23569 42820 23581 42823
rect 23348 42792 23581 42820
rect 23348 42780 23354 42792
rect 23569 42789 23581 42792
rect 23615 42789 23627 42823
rect 23569 42783 23627 42789
rect 23658 42780 23664 42832
rect 23716 42820 23722 42832
rect 24946 42820 24952 42832
rect 23716 42792 24952 42820
rect 23716 42780 23722 42792
rect 24946 42780 24952 42792
rect 25004 42780 25010 42832
rect 35894 42780 35900 42832
rect 35952 42820 35958 42832
rect 41598 42820 41604 42832
rect 35952 42792 41604 42820
rect 35952 42780 35958 42792
rect 41598 42780 41604 42792
rect 41656 42780 41662 42832
rect 41782 42780 41788 42832
rect 41840 42820 41846 42832
rect 41877 42823 41935 42829
rect 41877 42820 41889 42823
rect 41840 42792 41889 42820
rect 41840 42780 41846 42792
rect 41877 42789 41889 42792
rect 41923 42789 41935 42823
rect 41877 42783 41935 42789
rect 20349 42755 20407 42761
rect 20349 42721 20361 42755
rect 20395 42721 20407 42755
rect 20622 42752 20628 42764
rect 20583 42724 20628 42752
rect 20349 42715 20407 42721
rect 20254 42684 20260 42696
rect 20215 42656 20260 42684
rect 20254 42644 20260 42656
rect 20312 42644 20318 42696
rect 20364 42684 20392 42715
rect 20622 42712 20628 42724
rect 20680 42712 20686 42764
rect 21008 42724 21312 42752
rect 21008 42684 21036 42724
rect 21174 42684 21180 42696
rect 20364 42656 21036 42684
rect 21135 42656 21180 42684
rect 21174 42644 21180 42656
rect 21232 42644 21238 42696
rect 21284 42684 21312 42724
rect 23382 42712 23388 42764
rect 23440 42752 23446 42764
rect 25317 42755 25375 42761
rect 25317 42752 25329 42755
rect 23440 42724 25329 42752
rect 23440 42712 23446 42724
rect 25317 42721 25329 42724
rect 25363 42721 25375 42755
rect 25317 42715 25375 42721
rect 30561 42755 30619 42761
rect 30561 42721 30573 42755
rect 30607 42752 30619 42755
rect 30926 42752 30932 42764
rect 30607 42724 30932 42752
rect 30607 42721 30619 42724
rect 30561 42715 30619 42721
rect 30926 42712 30932 42724
rect 30984 42752 30990 42764
rect 31938 42752 31944 42764
rect 30984 42724 31800 42752
rect 31899 42724 31944 42752
rect 30984 42712 30990 42724
rect 22830 42684 22836 42696
rect 21284 42656 22836 42684
rect 22830 42644 22836 42656
rect 22888 42644 22894 42696
rect 23474 42684 23480 42696
rect 23435 42656 23480 42684
rect 23474 42644 23480 42656
rect 23532 42644 23538 42696
rect 23750 42644 23756 42696
rect 23808 42684 23814 42696
rect 24302 42684 24308 42696
rect 23808 42656 24308 42684
rect 23808 42644 23814 42656
rect 24302 42644 24308 42656
rect 24360 42644 24366 42696
rect 24397 42687 24455 42693
rect 24397 42653 24409 42687
rect 24443 42684 24455 42687
rect 24486 42684 24492 42696
rect 24443 42656 24492 42684
rect 24443 42653 24455 42656
rect 24397 42647 24455 42653
rect 21266 42576 21272 42628
rect 21324 42616 21330 42628
rect 21422 42619 21480 42625
rect 21422 42616 21434 42619
rect 21324 42588 21434 42616
rect 21324 42576 21330 42588
rect 21422 42585 21434 42588
rect 21468 42585 21480 42619
rect 21422 42579 21480 42585
rect 23293 42619 23351 42625
rect 23293 42585 23305 42619
rect 23339 42616 23351 42619
rect 24412 42616 24440 42647
rect 24486 42644 24492 42656
rect 24544 42644 24550 42696
rect 24670 42684 24676 42696
rect 24631 42656 24676 42684
rect 24670 42644 24676 42656
rect 24728 42644 24734 42696
rect 28074 42644 28080 42696
rect 28132 42684 28138 42696
rect 28261 42687 28319 42693
rect 28261 42684 28273 42687
rect 28132 42656 28273 42684
rect 28132 42644 28138 42656
rect 28261 42653 28273 42656
rect 28307 42653 28319 42687
rect 28261 42647 28319 42653
rect 28994 42644 29000 42696
rect 29052 42684 29058 42696
rect 29733 42687 29791 42693
rect 29733 42684 29745 42687
rect 29052 42656 29745 42684
rect 29052 42644 29058 42656
rect 29733 42653 29745 42656
rect 29779 42653 29791 42687
rect 30190 42684 30196 42696
rect 30151 42656 30196 42684
rect 29733 42647 29791 42653
rect 30190 42644 30196 42656
rect 30248 42644 30254 42696
rect 30377 42687 30435 42693
rect 30377 42653 30389 42687
rect 30423 42684 30435 42687
rect 31294 42684 31300 42696
rect 30423 42656 31300 42684
rect 30423 42653 30435 42656
rect 30377 42647 30435 42653
rect 31294 42644 31300 42656
rect 31352 42644 31358 42696
rect 31570 42684 31576 42696
rect 31531 42656 31576 42684
rect 31570 42644 31576 42656
rect 31628 42644 31634 42696
rect 31772 42693 31800 42724
rect 31938 42712 31944 42724
rect 31996 42712 32002 42764
rect 32674 42752 32680 42764
rect 32635 42724 32680 42752
rect 32674 42712 32680 42724
rect 32732 42712 32738 42764
rect 37550 42752 37556 42764
rect 37511 42724 37556 42752
rect 37550 42712 37556 42724
rect 37608 42712 37614 42764
rect 38378 42752 38384 42764
rect 38339 42724 38384 42752
rect 38378 42712 38384 42724
rect 38436 42712 38442 42764
rect 41984 42761 42012 42860
rect 42242 42848 42248 42860
rect 42300 42848 42306 42900
rect 42613 42891 42671 42897
rect 42613 42857 42625 42891
rect 42659 42857 42671 42891
rect 42613 42851 42671 42857
rect 42628 42820 42656 42851
rect 42702 42848 42708 42900
rect 42760 42888 42766 42900
rect 45370 42888 45376 42900
rect 42760 42860 45376 42888
rect 42760 42848 42766 42860
rect 45370 42848 45376 42860
rect 45428 42888 45434 42900
rect 46382 42888 46388 42900
rect 45428 42860 46388 42888
rect 45428 42848 45434 42860
rect 46382 42848 46388 42860
rect 46440 42848 46446 42900
rect 46661 42891 46719 42897
rect 46661 42857 46673 42891
rect 46707 42888 46719 42891
rect 46750 42888 46756 42900
rect 46707 42860 46756 42888
rect 46707 42857 46719 42860
rect 46661 42851 46719 42857
rect 46750 42848 46756 42860
rect 46808 42848 46814 42900
rect 48225 42891 48283 42897
rect 48225 42857 48237 42891
rect 48271 42888 48283 42891
rect 49786 42888 49792 42900
rect 48271 42860 49792 42888
rect 48271 42857 48283 42860
rect 48225 42851 48283 42857
rect 49786 42848 49792 42860
rect 49844 42848 49850 42900
rect 51353 42891 51411 42897
rect 51353 42857 51365 42891
rect 51399 42888 51411 42891
rect 51442 42888 51448 42900
rect 51399 42860 51448 42888
rect 51399 42857 51411 42860
rect 51353 42851 51411 42857
rect 51442 42848 51448 42860
rect 51500 42848 51506 42900
rect 52914 42848 52920 42900
rect 52972 42888 52978 42900
rect 53101 42891 53159 42897
rect 53101 42888 53113 42891
rect 52972 42860 53113 42888
rect 52972 42848 52978 42860
rect 53101 42857 53113 42860
rect 53147 42857 53159 42891
rect 55398 42888 55404 42900
rect 55359 42860 55404 42888
rect 53101 42851 53159 42857
rect 55398 42848 55404 42860
rect 55456 42848 55462 42900
rect 42628 42792 42840 42820
rect 42812 42764 42840 42792
rect 44266 42780 44272 42832
rect 44324 42820 44330 42832
rect 54754 42820 54760 42832
rect 44324 42792 54760 42820
rect 44324 42780 44330 42792
rect 54754 42780 54760 42792
rect 54812 42780 54818 42832
rect 41969 42755 42027 42761
rect 41969 42721 41981 42755
rect 42015 42721 42027 42755
rect 41969 42715 42027 42721
rect 42794 42712 42800 42764
rect 42852 42712 42858 42764
rect 44450 42712 44456 42764
rect 44508 42752 44514 42764
rect 45741 42755 45799 42761
rect 45741 42752 45753 42755
rect 44508 42724 45753 42752
rect 44508 42712 44514 42724
rect 45741 42721 45753 42724
rect 45787 42721 45799 42755
rect 47213 42755 47271 42761
rect 47213 42752 47225 42755
rect 45741 42715 45799 42721
rect 46584 42724 47225 42752
rect 46584 42696 46612 42724
rect 47213 42721 47225 42724
rect 47259 42721 47271 42755
rect 47213 42715 47271 42721
rect 52825 42755 52883 42761
rect 52825 42721 52837 42755
rect 52871 42721 52883 42755
rect 52825 42715 52883 42721
rect 31757 42687 31815 42693
rect 31757 42653 31769 42687
rect 31803 42684 31815 42687
rect 32493 42687 32551 42693
rect 32493 42684 32505 42687
rect 31803 42656 32505 42684
rect 31803 42653 31815 42656
rect 31757 42647 31815 42653
rect 32493 42653 32505 42656
rect 32539 42653 32551 42687
rect 34698 42684 34704 42696
rect 34659 42656 34704 42684
rect 32493 42647 32551 42653
rect 34698 42644 34704 42656
rect 34756 42644 34762 42696
rect 34968 42687 35026 42693
rect 34968 42653 34980 42687
rect 35014 42684 35026 42687
rect 36722 42684 36728 42696
rect 35014 42656 36728 42684
rect 35014 42653 35026 42656
rect 34968 42647 35026 42653
rect 36722 42644 36728 42656
rect 36780 42644 36786 42696
rect 37461 42687 37519 42693
rect 37461 42653 37473 42687
rect 37507 42653 37519 42687
rect 37461 42647 37519 42653
rect 38473 42687 38531 42693
rect 38473 42653 38485 42687
rect 38519 42684 38531 42687
rect 38562 42684 38568 42696
rect 38519 42656 38568 42684
rect 38519 42653 38531 42656
rect 38473 42647 38531 42653
rect 23339 42588 24440 42616
rect 25584 42619 25642 42625
rect 23339 42585 23351 42588
rect 23293 42579 23351 42585
rect 25584 42585 25596 42619
rect 25630 42616 25642 42619
rect 25774 42616 25780 42628
rect 25630 42588 25780 42616
rect 25630 42585 25642 42588
rect 25584 42579 25642 42585
rect 25774 42576 25780 42588
rect 25832 42576 25838 42628
rect 27249 42619 27307 42625
rect 27249 42585 27261 42619
rect 27295 42585 27307 42619
rect 27249 42579 27307 42585
rect 24486 42548 24492 42560
rect 24544 42557 24550 42560
rect 24453 42520 24492 42548
rect 24486 42508 24492 42520
rect 24544 42511 24553 42557
rect 24581 42551 24639 42557
rect 24581 42517 24593 42551
rect 24627 42548 24639 42551
rect 26697 42551 26755 42557
rect 26697 42548 26709 42551
rect 24627 42520 26709 42548
rect 24627 42517 24639 42520
rect 24581 42511 24639 42517
rect 26697 42517 26709 42520
rect 26743 42548 26755 42551
rect 27264 42548 27292 42579
rect 27430 42576 27436 42628
rect 27488 42616 27494 42628
rect 27488 42588 31754 42616
rect 27488 42576 27494 42588
rect 26743 42520 27292 42548
rect 28077 42551 28135 42557
rect 26743 42517 26755 42520
rect 26697 42511 26755 42517
rect 28077 42517 28089 42551
rect 28123 42548 28135 42551
rect 29362 42548 29368 42560
rect 28123 42520 29368 42548
rect 28123 42517 28135 42520
rect 28077 42511 28135 42517
rect 24544 42508 24550 42511
rect 29362 42508 29368 42520
rect 29420 42508 29426 42560
rect 29454 42508 29460 42560
rect 29512 42548 29518 42560
rect 29549 42551 29607 42557
rect 29549 42548 29561 42551
rect 29512 42520 29561 42548
rect 29512 42508 29518 42520
rect 29549 42517 29561 42520
rect 29595 42517 29607 42551
rect 31726 42548 31754 42588
rect 32306 42548 32312 42560
rect 31726 42520 32312 42548
rect 29549 42511 29607 42517
rect 32306 42508 32312 42520
rect 32364 42548 32370 42560
rect 32950 42548 32956 42560
rect 32364 42520 32956 42548
rect 32364 42508 32370 42520
rect 32950 42508 32956 42520
rect 33008 42508 33014 42560
rect 36078 42548 36084 42560
rect 36039 42520 36084 42548
rect 36078 42508 36084 42520
rect 36136 42508 36142 42560
rect 37476 42548 37504 42647
rect 38562 42644 38568 42656
rect 38620 42644 38626 42696
rect 41414 42644 41420 42696
rect 41472 42693 41478 42696
rect 41472 42687 41508 42693
rect 41496 42653 41508 42687
rect 41472 42647 41508 42653
rect 41472 42644 41478 42647
rect 42058 42644 42064 42696
rect 42116 42684 42122 42696
rect 42429 42687 42487 42693
rect 42429 42684 42441 42687
rect 42116 42656 42441 42684
rect 42116 42644 42122 42656
rect 42429 42653 42441 42656
rect 42475 42653 42487 42687
rect 42429 42647 42487 42653
rect 42613 42687 42671 42693
rect 42613 42653 42625 42687
rect 42659 42684 42671 42687
rect 44358 42684 44364 42696
rect 42659 42656 44364 42684
rect 42659 42653 42671 42656
rect 42613 42647 42671 42653
rect 44358 42644 44364 42656
rect 44416 42644 44422 42696
rect 45002 42684 45008 42696
rect 44963 42656 45008 42684
rect 45002 42644 45008 42656
rect 45060 42644 45066 42696
rect 45186 42684 45192 42696
rect 45099 42656 45192 42684
rect 45186 42644 45192 42656
rect 45244 42644 45250 42696
rect 45281 42687 45339 42693
rect 45281 42653 45293 42687
rect 45327 42653 45339 42687
rect 45281 42647 45339 42653
rect 38654 42616 38660 42628
rect 38567 42588 38660 42616
rect 38626 42576 38660 42588
rect 38712 42616 38718 42628
rect 39666 42616 39672 42628
rect 38712 42588 39672 42616
rect 38712 42576 38718 42588
rect 39666 42576 39672 42588
rect 39724 42576 39730 42628
rect 43070 42576 43076 42628
rect 43128 42616 43134 42628
rect 45204 42616 45232 42644
rect 43128 42588 45232 42616
rect 43128 42576 43134 42588
rect 38626 42548 38654 42576
rect 37476 42520 38654 42548
rect 41138 42508 41144 42560
rect 41196 42548 41202 42560
rect 41509 42551 41567 42557
rect 41509 42548 41521 42551
rect 41196 42520 41521 42548
rect 41196 42508 41202 42520
rect 41509 42517 41521 42520
rect 41555 42517 41567 42551
rect 41509 42511 41567 42517
rect 42797 42551 42855 42557
rect 42797 42517 42809 42551
rect 42843 42548 42855 42551
rect 42886 42548 42892 42560
rect 42843 42520 42892 42548
rect 42843 42517 42855 42520
rect 42797 42511 42855 42517
rect 42886 42508 42892 42520
rect 42944 42508 42950 42560
rect 45186 42508 45192 42560
rect 45244 42548 45250 42560
rect 45296 42548 45324 42647
rect 45370 42644 45376 42696
rect 45428 42684 45434 42696
rect 45554 42684 45560 42696
rect 45428 42656 45473 42684
rect 45515 42656 45560 42684
rect 45428 42644 45434 42656
rect 45554 42644 45560 42656
rect 45612 42644 45618 42696
rect 46293 42687 46351 42693
rect 46293 42653 46305 42687
rect 46339 42684 46351 42687
rect 46566 42684 46572 42696
rect 46339 42656 46572 42684
rect 46339 42653 46351 42656
rect 46293 42647 46351 42653
rect 46566 42644 46572 42656
rect 46624 42644 46630 42696
rect 47118 42684 47124 42696
rect 47079 42656 47124 42684
rect 47118 42644 47124 42656
rect 47176 42644 47182 42696
rect 47302 42684 47308 42696
rect 47263 42656 47308 42684
rect 47302 42644 47308 42656
rect 47360 42644 47366 42696
rect 48130 42684 48136 42696
rect 48091 42656 48136 42684
rect 48130 42644 48136 42656
rect 48188 42644 48194 42696
rect 48314 42684 48320 42696
rect 48275 42656 48320 42684
rect 48314 42644 48320 42656
rect 48372 42644 48378 42696
rect 49970 42644 49976 42696
rect 50028 42684 50034 42696
rect 51261 42687 51319 42693
rect 51261 42684 51273 42687
rect 50028 42656 51273 42684
rect 50028 42644 50034 42656
rect 51261 42653 51273 42656
rect 51307 42653 51319 42687
rect 51261 42647 51319 42653
rect 51445 42687 51503 42693
rect 51445 42653 51457 42687
rect 51491 42653 51503 42687
rect 51445 42647 51503 42653
rect 52733 42687 52791 42693
rect 52733 42653 52745 42687
rect 52779 42653 52791 42687
rect 52840 42684 52868 42715
rect 53834 42712 53840 42764
rect 53892 42752 53898 42764
rect 54389 42755 54447 42761
rect 54389 42752 54401 42755
rect 53892 42724 54401 42752
rect 53892 42712 53898 42724
rect 54389 42721 54401 42724
rect 54435 42721 54447 42755
rect 54389 42715 54447 42721
rect 56505 42755 56563 42761
rect 56505 42721 56517 42755
rect 56551 42752 56563 42755
rect 56870 42752 56876 42764
rect 56551 42724 56876 42752
rect 56551 42721 56563 42724
rect 56505 42715 56563 42721
rect 56870 42712 56876 42724
rect 56928 42712 56934 42764
rect 57882 42752 57888 42764
rect 57843 42724 57888 42752
rect 57882 42712 57888 42724
rect 57940 42712 57946 42764
rect 53466 42684 53472 42696
rect 52840 42656 53472 42684
rect 52733 42647 52791 42653
rect 46474 42616 46480 42628
rect 46435 42588 46480 42616
rect 46474 42576 46480 42588
rect 46532 42576 46538 42628
rect 48332 42616 48360 42644
rect 50614 42616 50620 42628
rect 46584 42588 48360 42616
rect 50575 42588 50620 42616
rect 46584 42548 46612 42588
rect 50614 42576 50620 42588
rect 50672 42576 50678 42628
rect 50798 42576 50804 42628
rect 50856 42616 50862 42628
rect 51460 42616 51488 42647
rect 50856 42588 51488 42616
rect 52748 42616 52776 42647
rect 53466 42644 53472 42656
rect 53524 42644 53530 42696
rect 55582 42684 55588 42696
rect 55543 42656 55588 42684
rect 55582 42644 55588 42656
rect 55640 42644 55646 42696
rect 56321 42687 56379 42693
rect 56321 42653 56333 42687
rect 56367 42653 56379 42687
rect 56321 42647 56379 42653
rect 53098 42616 53104 42628
rect 52748 42588 53104 42616
rect 50856 42576 50862 42588
rect 53098 42576 53104 42588
rect 53156 42576 53162 42628
rect 54018 42616 54024 42628
rect 53979 42588 54024 42616
rect 54018 42576 54024 42588
rect 54076 42576 54082 42628
rect 54205 42619 54263 42625
rect 54205 42585 54217 42619
rect 54251 42616 54263 42619
rect 54386 42616 54392 42628
rect 54251 42588 54392 42616
rect 54251 42585 54263 42588
rect 54205 42579 54263 42585
rect 45244 42520 46612 42548
rect 45244 42508 45250 42520
rect 48222 42508 48228 42560
rect 48280 42548 48286 42560
rect 50709 42551 50767 42557
rect 50709 42548 50721 42551
rect 48280 42520 50721 42548
rect 48280 42508 48286 42520
rect 50709 42517 50721 42520
rect 50755 42517 50767 42551
rect 50709 42511 50767 42517
rect 51534 42508 51540 42560
rect 51592 42548 51598 42560
rect 54220 42548 54248 42579
rect 54386 42576 54392 42588
rect 54444 42576 54450 42628
rect 55306 42616 55312 42628
rect 55267 42588 55312 42616
rect 55306 42576 55312 42588
rect 55364 42576 55370 42628
rect 55490 42616 55496 42628
rect 55451 42588 55496 42616
rect 55490 42576 55496 42588
rect 55548 42576 55554 42628
rect 56336 42616 56364 42647
rect 58066 42616 58072 42628
rect 56336 42588 58072 42616
rect 58066 42576 58072 42588
rect 58124 42576 58130 42628
rect 51592 42520 54248 42548
rect 51592 42508 51598 42520
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 20254 42304 20260 42356
rect 20312 42344 20318 42356
rect 20901 42347 20959 42353
rect 20901 42344 20913 42347
rect 20312 42316 20913 42344
rect 20312 42304 20318 42316
rect 20901 42313 20913 42316
rect 20947 42344 20959 42347
rect 23474 42344 23480 42356
rect 20947 42316 23480 42344
rect 20947 42313 20959 42316
rect 20901 42307 20959 42313
rect 23474 42304 23480 42316
rect 23532 42304 23538 42356
rect 25222 42344 25228 42356
rect 25183 42316 25228 42344
rect 25222 42304 25228 42316
rect 25280 42304 25286 42356
rect 25774 42344 25780 42356
rect 25735 42316 25780 42344
rect 25774 42304 25780 42316
rect 25832 42304 25838 42356
rect 29546 42344 29552 42356
rect 29507 42316 29552 42344
rect 29546 42304 29552 42316
rect 29604 42304 29610 42356
rect 32674 42344 32680 42356
rect 32232 42316 32680 42344
rect 21174 42276 21180 42288
rect 19536 42248 21180 42276
rect 19536 42217 19564 42248
rect 21174 42236 21180 42248
rect 21232 42276 21238 42288
rect 22370 42276 22376 42288
rect 21232 42248 22376 42276
rect 21232 42236 21238 42248
rect 22370 42236 22376 42248
rect 22428 42276 22434 42288
rect 23382 42276 23388 42288
rect 22428 42248 23388 42276
rect 22428 42236 22434 42248
rect 23382 42236 23388 42248
rect 23440 42276 23446 42288
rect 23440 42248 23888 42276
rect 23440 42236 23446 42248
rect 19521 42211 19579 42217
rect 19521 42177 19533 42211
rect 19567 42177 19579 42211
rect 19521 42171 19579 42177
rect 19788 42211 19846 42217
rect 19788 42177 19800 42211
rect 19834 42208 19846 42211
rect 20162 42208 20168 42220
rect 19834 42180 20168 42208
rect 19834 42177 19846 42180
rect 19788 42171 19846 42177
rect 20162 42168 20168 42180
rect 20220 42168 20226 42220
rect 22002 42208 22008 42220
rect 21963 42180 22008 42208
rect 22002 42168 22008 42180
rect 22060 42168 22066 42220
rect 23860 42217 23888 42248
rect 23845 42211 23903 42217
rect 23845 42177 23857 42211
rect 23891 42177 23903 42211
rect 23845 42171 23903 42177
rect 23934 42168 23940 42220
rect 23992 42208 23998 42220
rect 24101 42211 24159 42217
rect 24101 42208 24113 42211
rect 23992 42180 24113 42208
rect 23992 42168 23998 42180
rect 24101 42177 24113 42180
rect 24147 42177 24159 42211
rect 25958 42208 25964 42220
rect 25919 42180 25964 42208
rect 24101 42171 24159 42177
rect 25958 42168 25964 42180
rect 26016 42168 26022 42220
rect 26234 42208 26240 42220
rect 26195 42180 26240 42208
rect 26234 42168 26240 42180
rect 26292 42168 26298 42220
rect 26326 42168 26332 42220
rect 26384 42208 26390 42220
rect 26421 42211 26479 42217
rect 26421 42208 26433 42211
rect 26384 42180 26433 42208
rect 26384 42168 26390 42180
rect 26421 42177 26433 42180
rect 26467 42208 26479 42211
rect 27430 42208 27436 42220
rect 26467 42180 27436 42208
rect 26467 42177 26479 42180
rect 26421 42171 26479 42177
rect 27430 42168 27436 42180
rect 27488 42168 27494 42220
rect 27522 42168 27528 42220
rect 27580 42208 27586 42220
rect 28258 42208 28264 42220
rect 27580 42180 27625 42208
rect 28219 42180 28264 42208
rect 27580 42168 27586 42180
rect 28258 42168 28264 42180
rect 28316 42168 28322 42220
rect 29822 42168 29828 42220
rect 29880 42208 29886 42220
rect 30653 42211 30711 42217
rect 30653 42208 30665 42211
rect 29880 42180 30665 42208
rect 29880 42168 29886 42180
rect 30653 42177 30665 42180
rect 30699 42177 30711 42211
rect 30653 42171 30711 42177
rect 31205 42211 31263 42217
rect 31205 42177 31217 42211
rect 31251 42177 31263 42211
rect 31386 42208 31392 42220
rect 31347 42180 31392 42208
rect 31205 42171 31263 42177
rect 20622 42100 20628 42152
rect 20680 42140 20686 42152
rect 21913 42143 21971 42149
rect 21913 42140 21925 42143
rect 20680 42112 21925 42140
rect 20680 42100 20686 42112
rect 21913 42109 21925 42112
rect 21959 42109 21971 42143
rect 21913 42103 21971 42109
rect 30466 42100 30472 42152
rect 30524 42140 30530 42152
rect 31220 42140 31248 42171
rect 31386 42168 31392 42180
rect 31444 42168 31450 42220
rect 32125 42211 32183 42217
rect 32125 42177 32137 42211
rect 32171 42177 32183 42211
rect 32232 42208 32260 42316
rect 32674 42304 32680 42316
rect 32732 42304 32738 42356
rect 35618 42344 35624 42356
rect 35579 42316 35624 42344
rect 35618 42304 35624 42316
rect 35676 42304 35682 42356
rect 38657 42347 38715 42353
rect 38657 42313 38669 42347
rect 38703 42344 38715 42347
rect 38930 42344 38936 42356
rect 38703 42316 38936 42344
rect 38703 42313 38715 42316
rect 38657 42307 38715 42313
rect 38930 42304 38936 42316
rect 38988 42304 38994 42356
rect 41699 42347 41757 42353
rect 41699 42344 41711 42347
rect 39316 42316 41711 42344
rect 39316 42288 39344 42316
rect 41699 42313 41711 42316
rect 41745 42344 41757 42347
rect 42058 42344 42064 42356
rect 41745 42316 42064 42344
rect 41745 42313 41757 42316
rect 41699 42307 41757 42313
rect 42058 42304 42064 42316
rect 42116 42304 42122 42356
rect 42794 42344 42800 42356
rect 42755 42316 42800 42344
rect 42794 42304 42800 42316
rect 42852 42304 42858 42356
rect 47118 42304 47124 42356
rect 47176 42344 47182 42356
rect 49234 42344 49240 42356
rect 47176 42316 49240 42344
rect 47176 42304 47182 42316
rect 49234 42304 49240 42316
rect 49292 42304 49298 42356
rect 50062 42344 50068 42356
rect 50023 42316 50068 42344
rect 50062 42304 50068 42316
rect 50120 42304 50126 42356
rect 51813 42347 51871 42353
rect 51813 42313 51825 42347
rect 51859 42344 51871 42347
rect 52270 42344 52276 42356
rect 51859 42316 52276 42344
rect 51859 42313 51871 42316
rect 51813 42307 51871 42313
rect 52270 42304 52276 42316
rect 52328 42304 52334 42356
rect 54018 42304 54024 42356
rect 54076 42344 54082 42356
rect 54481 42347 54539 42353
rect 54481 42344 54493 42347
rect 54076 42316 54493 42344
rect 54076 42304 54082 42316
rect 54481 42313 54493 42316
rect 54527 42313 54539 42347
rect 54481 42307 54539 42313
rect 55401 42347 55459 42353
rect 55401 42313 55413 42347
rect 55447 42344 55459 42347
rect 55582 42344 55588 42356
rect 55447 42316 55588 42344
rect 55447 42313 55459 42316
rect 55401 42307 55459 42313
rect 55582 42304 55588 42316
rect 55640 42304 55646 42356
rect 56962 42344 56968 42356
rect 56923 42316 56968 42344
rect 56962 42304 56968 42316
rect 57020 42304 57026 42356
rect 32398 42276 32404 42288
rect 32359 42248 32404 42276
rect 32398 42236 32404 42248
rect 32456 42236 32462 42288
rect 34698 42276 34704 42288
rect 34256 42248 34704 42276
rect 32309 42211 32367 42217
rect 32309 42208 32321 42211
rect 32232 42180 32321 42208
rect 32125 42171 32183 42177
rect 32309 42177 32321 42180
rect 32355 42177 32367 42211
rect 32490 42208 32496 42220
rect 32451 42180 32496 42208
rect 32309 42171 32367 42177
rect 30524 42112 31248 42140
rect 32140 42140 32168 42171
rect 32490 42168 32496 42180
rect 32548 42168 32554 42220
rect 34256 42217 34284 42248
rect 34698 42236 34704 42248
rect 34756 42236 34762 42288
rect 39298 42276 39304 42288
rect 39211 42248 39304 42276
rect 39298 42236 39304 42248
rect 39356 42236 39362 42288
rect 41601 42279 41659 42285
rect 41601 42245 41613 42279
rect 41647 42276 41659 42279
rect 42426 42276 42432 42288
rect 41647 42248 42432 42276
rect 41647 42245 41659 42248
rect 41601 42239 41659 42245
rect 42426 42236 42432 42248
rect 42484 42236 42490 42288
rect 48590 42276 48596 42288
rect 42659 42245 42717 42251
rect 48551 42248 48596 42276
rect 42659 42242 42671 42245
rect 34241 42211 34299 42217
rect 34241 42177 34253 42211
rect 34287 42177 34299 42211
rect 34241 42171 34299 42177
rect 34508 42211 34566 42217
rect 34508 42177 34520 42211
rect 34554 42208 34566 42211
rect 35526 42208 35532 42220
rect 34554 42180 35532 42208
rect 34554 42177 34566 42180
rect 34508 42171 34566 42177
rect 35526 42168 35532 42180
rect 35584 42168 35590 42220
rect 37826 42168 37832 42220
rect 37884 42208 37890 42220
rect 38194 42208 38200 42220
rect 37884 42180 38200 42208
rect 37884 42168 37890 42180
rect 38194 42168 38200 42180
rect 38252 42208 38258 42220
rect 38289 42211 38347 42217
rect 38289 42208 38301 42211
rect 38252 42180 38301 42208
rect 38252 42168 38258 42180
rect 38289 42177 38301 42180
rect 38335 42177 38347 42211
rect 39114 42208 39120 42220
rect 39075 42180 39120 42208
rect 38289 42171 38347 42177
rect 39114 42168 39120 42180
rect 39172 42168 39178 42220
rect 40497 42211 40555 42217
rect 40497 42177 40509 42211
rect 40543 42177 40555 42211
rect 40497 42171 40555 42177
rect 40681 42211 40739 42217
rect 40681 42177 40693 42211
rect 40727 42208 40739 42211
rect 41138 42208 41144 42220
rect 40727 42180 41144 42208
rect 40727 42177 40739 42180
rect 40681 42171 40739 42177
rect 33502 42140 33508 42152
rect 32140 42112 33508 42140
rect 30524 42100 30530 42112
rect 33502 42100 33508 42112
rect 33560 42100 33566 42152
rect 38381 42143 38439 42149
rect 38381 42109 38393 42143
rect 38427 42140 38439 42143
rect 39485 42143 39543 42149
rect 39485 42140 39497 42143
rect 38427 42112 39497 42140
rect 38427 42109 38439 42112
rect 38381 42103 38439 42109
rect 39485 42109 39497 42112
rect 39531 42109 39543 42143
rect 40512 42140 40540 42171
rect 41138 42168 41144 42180
rect 41196 42168 41202 42220
rect 41785 42211 41843 42217
rect 41785 42177 41797 42211
rect 41831 42177 41843 42211
rect 41785 42171 41843 42177
rect 41690 42140 41696 42152
rect 40512 42112 41696 42140
rect 39485 42103 39543 42109
rect 41690 42100 41696 42112
rect 41748 42100 41754 42152
rect 32030 42032 32036 42084
rect 32088 42072 32094 42084
rect 32677 42075 32735 42081
rect 32677 42072 32689 42075
rect 32088 42044 32689 42072
rect 32088 42032 32094 42044
rect 32677 42041 32689 42044
rect 32723 42041 32735 42075
rect 32677 42035 32735 42041
rect 22278 42004 22284 42016
rect 22239 41976 22284 42004
rect 22278 41964 22284 41976
rect 22336 41964 22342 42016
rect 24578 41964 24584 42016
rect 24636 42004 24642 42016
rect 27706 42004 27712 42016
rect 24636 41976 27712 42004
rect 24636 41964 24642 41976
rect 27706 41964 27712 41976
rect 27764 41964 27770 42016
rect 30374 41964 30380 42016
rect 30432 42004 30438 42016
rect 30469 42007 30527 42013
rect 30469 42004 30481 42007
rect 30432 41976 30481 42004
rect 30432 41964 30438 41976
rect 30469 41973 30481 41976
rect 30515 41973 30527 42007
rect 31202 42004 31208 42016
rect 31163 41976 31208 42004
rect 30469 41967 30527 41973
rect 31202 41964 31208 41976
rect 31260 41964 31266 42016
rect 32398 41964 32404 42016
rect 32456 42004 32462 42016
rect 32766 42004 32772 42016
rect 32456 41976 32772 42004
rect 32456 41964 32462 41976
rect 32766 41964 32772 41976
rect 32824 41964 32830 42016
rect 39666 41964 39672 42016
rect 39724 42004 39730 42016
rect 40773 42007 40831 42013
rect 40773 42004 40785 42007
rect 39724 41976 40785 42004
rect 39724 41964 39730 41976
rect 40773 41973 40785 41976
rect 40819 41973 40831 42007
rect 41800 42004 41828 42171
rect 41874 42168 41880 42220
rect 41932 42208 41938 42220
rect 42644 42211 42671 42242
rect 42705 42211 42717 42245
rect 48590 42236 48596 42248
rect 48648 42236 48654 42288
rect 56502 42236 56508 42288
rect 56560 42276 56566 42288
rect 56560 42248 57100 42276
rect 56560 42236 56566 42248
rect 42644 42208 42717 42211
rect 43254 42208 43260 42220
rect 41932 42205 42717 42208
rect 41932 42180 42672 42205
rect 43215 42180 43260 42208
rect 41932 42168 41938 42180
rect 43254 42168 43260 42180
rect 43312 42168 43318 42220
rect 43438 42208 43444 42220
rect 43399 42180 43444 42208
rect 43438 42168 43444 42180
rect 43496 42168 43502 42220
rect 47762 42208 47768 42220
rect 47723 42180 47768 42208
rect 47762 42168 47768 42180
rect 47820 42168 47826 42220
rect 47857 42211 47915 42217
rect 47857 42177 47869 42211
rect 47903 42208 47915 42211
rect 48498 42208 48504 42220
rect 47903 42180 48504 42208
rect 47903 42177 47915 42180
rect 47857 42171 47915 42177
rect 48498 42168 48504 42180
rect 48556 42168 48562 42220
rect 46474 42100 46480 42152
rect 46532 42140 46538 42152
rect 48608 42140 48636 42236
rect 48685 42211 48743 42217
rect 48685 42177 48697 42211
rect 48731 42208 48743 42211
rect 48866 42208 48872 42220
rect 48731 42180 48872 42208
rect 48731 42177 48743 42180
rect 48685 42171 48743 42177
rect 48866 42168 48872 42180
rect 48924 42168 48930 42220
rect 49970 42208 49976 42220
rect 49931 42180 49976 42208
rect 49970 42168 49976 42180
rect 50028 42168 50034 42220
rect 50157 42211 50215 42217
rect 50157 42177 50169 42211
rect 50203 42208 50215 42211
rect 50798 42208 50804 42220
rect 50203 42180 50804 42208
rect 50203 42177 50215 42180
rect 50157 42171 50215 42177
rect 46532 42112 48636 42140
rect 46532 42100 46538 42112
rect 49786 42100 49792 42152
rect 49844 42140 49850 42152
rect 50172 42140 50200 42171
rect 50798 42168 50804 42180
rect 50856 42168 50862 42220
rect 51534 42168 51540 42220
rect 51592 42208 51598 42220
rect 51721 42211 51779 42217
rect 51721 42208 51733 42211
rect 51592 42180 51733 42208
rect 51592 42168 51598 42180
rect 51721 42177 51733 42180
rect 51767 42177 51779 42211
rect 51902 42208 51908 42220
rect 51863 42180 51908 42208
rect 51721 42171 51779 42177
rect 51902 42168 51908 42180
rect 51960 42168 51966 42220
rect 54110 42208 54116 42220
rect 54071 42180 54116 42208
rect 54110 42168 54116 42180
rect 54168 42168 54174 42220
rect 54941 42211 54999 42217
rect 54941 42208 54953 42211
rect 54220 42180 54953 42208
rect 54220 42149 54248 42180
rect 54941 42177 54953 42180
rect 54987 42208 54999 42211
rect 55122 42208 55128 42220
rect 54987 42180 55128 42208
rect 54987 42177 54999 42180
rect 54941 42171 54999 42177
rect 55122 42168 55128 42180
rect 55180 42168 55186 42220
rect 57072 42217 57100 42248
rect 56873 42211 56931 42217
rect 56873 42177 56885 42211
rect 56919 42177 56931 42211
rect 56873 42171 56931 42177
rect 57057 42211 57115 42217
rect 57057 42177 57069 42211
rect 57103 42177 57115 42211
rect 58066 42208 58072 42220
rect 58027 42180 58072 42208
rect 57057 42171 57115 42177
rect 49844 42112 50200 42140
rect 54205 42143 54263 42149
rect 49844 42100 49850 42112
rect 54205 42109 54217 42143
rect 54251 42109 54263 42143
rect 56888 42140 56916 42171
rect 58066 42168 58072 42180
rect 58124 42168 58130 42220
rect 57330 42140 57336 42152
rect 56888 42112 57336 42140
rect 54205 42103 54263 42109
rect 57330 42100 57336 42112
rect 57388 42100 57394 42152
rect 42426 42032 42432 42084
rect 42484 42072 42490 42084
rect 43257 42075 43315 42081
rect 43257 42072 43269 42075
rect 42484 42044 43269 42072
rect 42484 42032 42490 42044
rect 43257 42041 43269 42044
rect 43303 42041 43315 42075
rect 43257 42035 43315 42041
rect 47302 42032 47308 42084
rect 47360 42072 47366 42084
rect 47854 42072 47860 42084
rect 47360 42044 47860 42072
rect 47360 42032 47366 42044
rect 47854 42032 47860 42044
rect 47912 42072 47918 42084
rect 48041 42075 48099 42081
rect 48041 42072 48053 42075
rect 47912 42044 48053 42072
rect 47912 42032 47918 42044
rect 48041 42041 48053 42044
rect 48087 42041 48099 42075
rect 48041 42035 48099 42041
rect 50154 42032 50160 42084
rect 50212 42072 50218 42084
rect 50798 42072 50804 42084
rect 50212 42044 50804 42072
rect 50212 42032 50218 42044
rect 50798 42032 50804 42044
rect 50856 42032 50862 42084
rect 42613 42007 42671 42013
rect 42613 42004 42625 42007
rect 41800 41976 42625 42004
rect 40773 41967 40831 41973
rect 42613 41973 42625 41976
rect 42659 42004 42671 42007
rect 42702 42004 42708 42016
rect 42659 41976 42708 42004
rect 42659 41973 42671 41976
rect 42613 41967 42671 41973
rect 42702 41964 42708 41976
rect 42760 41964 42766 42016
rect 54110 41964 54116 42016
rect 54168 42004 54174 42016
rect 55033 42007 55091 42013
rect 55033 42004 55045 42007
rect 54168 41976 55045 42004
rect 54168 41964 54174 41976
rect 55033 41973 55045 41976
rect 55079 41973 55091 42007
rect 55033 41967 55091 41973
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 20162 41800 20168 41812
rect 20123 41772 20168 41800
rect 20162 41760 20168 41772
rect 20220 41760 20226 41812
rect 20990 41800 20996 41812
rect 20456 41772 20996 41800
rect 20456 41732 20484 41772
rect 20990 41760 20996 41772
rect 21048 41760 21054 41812
rect 21266 41800 21272 41812
rect 21227 41772 21272 41800
rect 21266 41760 21272 41772
rect 21324 41760 21330 41812
rect 22002 41760 22008 41812
rect 22060 41800 22066 41812
rect 22373 41803 22431 41809
rect 22373 41800 22385 41803
rect 22060 41772 22385 41800
rect 22060 41760 22066 41772
rect 22373 41769 22385 41772
rect 22419 41769 22431 41803
rect 22373 41763 22431 41769
rect 23569 41803 23627 41809
rect 23569 41769 23581 41803
rect 23615 41800 23627 41803
rect 23934 41800 23940 41812
rect 23615 41772 23940 41800
rect 23615 41769 23627 41772
rect 23569 41763 23627 41769
rect 23934 41760 23940 41772
rect 23992 41760 23998 41812
rect 24946 41800 24952 41812
rect 24859 41772 24952 41800
rect 24946 41760 24952 41772
rect 25004 41800 25010 41812
rect 27522 41800 27528 41812
rect 25004 41772 27528 41800
rect 25004 41760 25010 41772
rect 27522 41760 27528 41772
rect 27580 41760 27586 41812
rect 28074 41800 28080 41812
rect 28035 41772 28080 41800
rect 28074 41760 28080 41772
rect 28132 41760 28138 41812
rect 28994 41800 29000 41812
rect 28955 41772 29000 41800
rect 28994 41760 29000 41772
rect 29052 41760 29058 41812
rect 31294 41760 31300 41812
rect 31352 41800 31358 41812
rect 31481 41803 31539 41809
rect 31481 41800 31493 41803
rect 31352 41772 31493 41800
rect 31352 41760 31358 41772
rect 31481 41769 31493 41772
rect 31527 41769 31539 41803
rect 33045 41803 33103 41809
rect 33045 41800 33057 41803
rect 31481 41763 31539 41769
rect 31588 41772 33057 41800
rect 19536 41704 20484 41732
rect 28905 41735 28963 41741
rect 19536 41605 19564 41704
rect 28905 41701 28917 41735
rect 28951 41732 28963 41735
rect 29914 41732 29920 41744
rect 28951 41704 29920 41732
rect 28951 41701 28963 41704
rect 28905 41695 28963 41701
rect 29914 41692 29920 41704
rect 29972 41692 29978 41744
rect 31202 41692 31208 41744
rect 31260 41732 31266 41744
rect 31588 41732 31616 41772
rect 33045 41769 33057 41772
rect 33091 41769 33103 41803
rect 33045 41763 33103 41769
rect 37093 41803 37151 41809
rect 37093 41769 37105 41803
rect 37139 41800 37151 41803
rect 38378 41800 38384 41812
rect 37139 41772 38384 41800
rect 37139 41769 37151 41772
rect 37093 41763 37151 41769
rect 38378 41760 38384 41772
rect 38436 41760 38442 41812
rect 42429 41803 42487 41809
rect 42429 41769 42441 41803
rect 42475 41800 42487 41803
rect 43254 41800 43260 41812
rect 42475 41772 43260 41800
rect 42475 41769 42487 41772
rect 42429 41763 42487 41769
rect 43254 41760 43260 41772
rect 43312 41760 43318 41812
rect 48314 41760 48320 41812
rect 48372 41800 48378 41812
rect 48593 41803 48651 41809
rect 48593 41800 48605 41803
rect 48372 41772 48605 41800
rect 48372 41760 48378 41772
rect 48593 41769 48605 41772
rect 48639 41769 48651 41803
rect 48593 41763 48651 41769
rect 56502 41760 56508 41812
rect 56560 41800 56566 41812
rect 56689 41803 56747 41809
rect 56689 41800 56701 41803
rect 56560 41772 56701 41800
rect 56560 41760 56566 41772
rect 56689 41769 56701 41772
rect 56735 41769 56747 41803
rect 56689 41763 56747 41769
rect 33594 41732 33600 41744
rect 31260 41704 31616 41732
rect 32140 41704 33600 41732
rect 31260 41692 31266 41704
rect 21174 41664 21180 41676
rect 20548 41636 21180 41664
rect 19521 41599 19579 41605
rect 19521 41565 19533 41599
rect 19567 41565 19579 41599
rect 19521 41559 19579 41565
rect 19705 41599 19763 41605
rect 19705 41565 19717 41599
rect 19751 41596 19763 41599
rect 19978 41596 19984 41608
rect 19751 41568 19984 41596
rect 19751 41565 19763 41568
rect 19705 41559 19763 41565
rect 19978 41556 19984 41568
rect 20036 41556 20042 41608
rect 20438 41596 20444 41608
rect 20399 41568 20444 41596
rect 20438 41556 20444 41568
rect 20496 41556 20502 41608
rect 20548 41605 20576 41636
rect 21174 41624 21180 41636
rect 21232 41664 21238 41676
rect 22370 41664 22376 41676
rect 21232 41636 21671 41664
rect 21232 41624 21238 41636
rect 20533 41599 20591 41605
rect 20533 41565 20545 41599
rect 20579 41565 20591 41599
rect 20533 41559 20591 41565
rect 20646 41599 20704 41605
rect 20646 41565 20658 41599
rect 20692 41596 20704 41599
rect 20692 41568 20760 41596
rect 20692 41565 20704 41568
rect 20646 41559 20704 41565
rect 20732 41528 20760 41568
rect 20806 41556 20812 41608
rect 20864 41596 20870 41608
rect 21643 41605 21671 41636
rect 21928 41636 22376 41664
rect 21928 41608 21956 41636
rect 22370 41624 22376 41636
rect 22428 41664 22434 41676
rect 25038 41664 25044 41676
rect 22428 41636 25044 41664
rect 22428 41624 22434 41636
rect 25038 41624 25044 41636
rect 25096 41624 25102 41676
rect 27709 41667 27767 41673
rect 27709 41633 27721 41667
rect 27755 41664 27767 41667
rect 27982 41664 27988 41676
rect 27755 41636 27988 41664
rect 27755 41633 27767 41636
rect 27709 41627 27767 41633
rect 21499 41599 21557 41605
rect 20864 41568 20909 41596
rect 20864 41556 20870 41568
rect 21499 41565 21511 41599
rect 21545 41565 21557 41599
rect 21499 41562 21557 41565
rect 21468 41559 21557 41562
rect 21634 41599 21692 41605
rect 21634 41565 21646 41599
rect 21680 41565 21692 41599
rect 21634 41559 21692 41565
rect 21468 41540 21542 41559
rect 21726 41556 21732 41608
rect 21784 41605 21790 41608
rect 21784 41596 21792 41605
rect 21784 41568 21829 41596
rect 21784 41559 21792 41568
rect 21784 41556 21790 41559
rect 21910 41556 21916 41608
rect 21968 41596 21974 41608
rect 21968 41568 22061 41596
rect 21968 41556 21974 41568
rect 22186 41556 22192 41608
rect 22244 41596 22250 41608
rect 22557 41599 22615 41605
rect 22557 41596 22569 41599
rect 22244 41568 22569 41596
rect 22244 41556 22250 41568
rect 22557 41565 22569 41568
rect 22603 41565 22615 41599
rect 22830 41596 22836 41608
rect 22791 41568 22836 41596
rect 22557 41559 22615 41565
rect 22830 41556 22836 41568
rect 22888 41556 22894 41608
rect 23845 41599 23903 41605
rect 23845 41565 23857 41599
rect 23891 41596 23903 41599
rect 24118 41596 24124 41608
rect 23891 41568 24124 41596
rect 23891 41565 23903 41568
rect 23845 41559 23903 41565
rect 24118 41556 24124 41568
rect 24176 41556 24182 41608
rect 24857 41599 24915 41605
rect 24857 41565 24869 41599
rect 24903 41596 24915 41599
rect 25222 41596 25228 41608
rect 24903 41568 25228 41596
rect 24903 41565 24915 41568
rect 24857 41559 24915 41565
rect 25222 41556 25228 41568
rect 25280 41556 25286 41608
rect 27065 41599 27123 41605
rect 27065 41565 27077 41599
rect 27111 41596 27123 41599
rect 27724 41596 27752 41627
rect 27982 41624 27988 41636
rect 28040 41624 28046 41676
rect 28534 41664 28540 41676
rect 28495 41636 28540 41664
rect 28534 41624 28540 41636
rect 28592 41624 28598 41676
rect 29362 41624 29368 41676
rect 29420 41664 29426 41676
rect 29420 41636 30236 41664
rect 29420 41624 29426 41636
rect 27111 41568 27752 41596
rect 27893 41599 27951 41605
rect 27111 41565 27123 41568
rect 27065 41559 27123 41565
rect 27893 41565 27905 41599
rect 27939 41596 27951 41599
rect 28902 41596 28908 41608
rect 27939 41568 28908 41596
rect 27939 41565 27951 41568
rect 27893 41559 27951 41565
rect 28902 41556 28908 41568
rect 28960 41556 28966 41608
rect 28994 41556 29000 41608
rect 29052 41596 29058 41608
rect 30101 41599 30159 41605
rect 30101 41596 30113 41599
rect 29052 41568 30113 41596
rect 29052 41556 29058 41568
rect 30101 41565 30113 41568
rect 30147 41565 30159 41599
rect 30208 41596 30236 41636
rect 32140 41605 32168 41704
rect 33594 41692 33600 41704
rect 33652 41692 33658 41744
rect 42518 41692 42524 41744
rect 42576 41732 42582 41744
rect 47857 41735 47915 41741
rect 42576 41704 47808 41732
rect 42576 41692 42582 41704
rect 32582 41664 32588 41676
rect 32543 41636 32588 41664
rect 32582 41624 32588 41636
rect 32640 41624 32646 41676
rect 38013 41667 38071 41673
rect 38013 41664 38025 41667
rect 37568 41636 38025 41664
rect 37568 41608 37596 41636
rect 38013 41633 38025 41636
rect 38059 41633 38071 41667
rect 45554 41664 45560 41676
rect 38013 41627 38071 41633
rect 45112 41636 45560 41664
rect 30357 41599 30415 41605
rect 30357 41596 30369 41599
rect 30208 41568 30369 41596
rect 30101 41559 30159 41565
rect 30357 41565 30369 41568
rect 30403 41565 30415 41599
rect 30357 41559 30415 41565
rect 32125 41599 32183 41605
rect 32125 41565 32137 41599
rect 32171 41565 32183 41599
rect 32310 41599 32368 41605
rect 32310 41586 32322 41599
rect 32356 41586 32368 41599
rect 32125 41559 32183 41565
rect 20732 41500 21220 41528
rect 19613 41463 19671 41469
rect 19613 41429 19625 41463
rect 19659 41460 19671 41463
rect 21082 41460 21088 41472
rect 19659 41432 21088 41460
rect 19659 41429 19671 41432
rect 19613 41423 19671 41429
rect 21082 41420 21088 41432
rect 21140 41420 21146 41472
rect 21192 41460 21220 41500
rect 21450 41488 21456 41540
rect 21508 41534 21542 41540
rect 21508 41488 21514 41534
rect 22738 41528 22744 41540
rect 22699 41500 22744 41528
rect 22738 41488 22744 41500
rect 22796 41488 22802 41540
rect 23569 41531 23627 41537
rect 23569 41497 23581 41531
rect 23615 41528 23627 41531
rect 24762 41528 24768 41540
rect 23615 41500 24768 41528
rect 23615 41497 23627 41500
rect 23569 41491 23627 41497
rect 24762 41488 24768 41500
rect 24820 41488 24826 41540
rect 31110 41488 31116 41540
rect 31168 41528 31174 41540
rect 31570 41528 31576 41540
rect 31168 41500 31576 41528
rect 31168 41488 31174 41500
rect 31570 41488 31576 41500
rect 31628 41528 31634 41540
rect 32217 41531 32275 41537
rect 32306 41534 32312 41586
rect 32364 41534 32370 41586
rect 32674 41556 32680 41608
rect 32732 41596 32738 41608
rect 33229 41599 33287 41605
rect 33229 41596 33241 41599
rect 32732 41568 33241 41596
rect 32732 41556 32738 41568
rect 33229 41565 33241 41568
rect 33275 41565 33287 41599
rect 33229 41559 33287 41565
rect 33505 41599 33563 41605
rect 33505 41565 33517 41599
rect 33551 41565 33563 41599
rect 37274 41596 37280 41608
rect 37235 41568 37280 41596
rect 33505 41559 33563 41565
rect 32217 41528 32229 41531
rect 31628 41500 32229 41528
rect 31628 41488 31634 41500
rect 32217 41497 32229 41500
rect 32263 41497 32275 41531
rect 32427 41531 32485 41537
rect 32427 41528 32439 41531
rect 32217 41491 32275 41497
rect 32416 41497 32439 41528
rect 32473 41497 32485 41531
rect 33520 41528 33548 41559
rect 37274 41556 37280 41568
rect 37332 41556 37338 41608
rect 37550 41596 37556 41608
rect 37511 41568 37556 41596
rect 37550 41556 37556 41568
rect 37608 41556 37614 41608
rect 37918 41556 37924 41608
rect 37976 41596 37982 41608
rect 38197 41599 38255 41605
rect 38197 41596 38209 41599
rect 37976 41568 38209 41596
rect 37976 41556 37982 41568
rect 38197 41565 38209 41568
rect 38243 41565 38255 41599
rect 38197 41559 38255 41565
rect 38473 41599 38531 41605
rect 38473 41565 38485 41599
rect 38519 41565 38531 41599
rect 38473 41559 38531 41565
rect 38657 41599 38715 41605
rect 38657 41565 38669 41599
rect 38703 41596 38715 41599
rect 39298 41596 39304 41608
rect 38703 41568 39304 41596
rect 38703 41565 38715 41568
rect 38657 41559 38715 41565
rect 32416 41491 32485 41497
rect 32600 41500 33548 41528
rect 38488 41528 38516 41559
rect 39298 41556 39304 41568
rect 39356 41556 39362 41608
rect 42426 41596 42432 41608
rect 42387 41568 42432 41596
rect 42426 41556 42432 41568
rect 42484 41556 42490 41608
rect 42613 41599 42671 41605
rect 42613 41565 42625 41599
rect 42659 41596 42671 41599
rect 43162 41596 43168 41608
rect 42659 41568 43168 41596
rect 42659 41565 42671 41568
rect 42613 41559 42671 41565
rect 43162 41556 43168 41568
rect 43220 41556 43226 41608
rect 45112 41605 45140 41636
rect 45554 41624 45560 41636
rect 45612 41664 45618 41676
rect 47670 41664 47676 41676
rect 45612 41636 47676 41664
rect 45612 41624 45618 41636
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 47780 41664 47808 41704
rect 47857 41701 47869 41735
rect 47903 41732 47915 41735
rect 47946 41732 47952 41744
rect 47903 41704 47952 41732
rect 47903 41701 47915 41704
rect 47857 41695 47915 41701
rect 47946 41692 47952 41704
rect 48004 41692 48010 41744
rect 51074 41664 51080 41676
rect 47780 41636 51080 41664
rect 51074 41624 51080 41636
rect 51132 41624 51138 41676
rect 45097 41599 45155 41605
rect 45097 41565 45109 41599
rect 45143 41565 45155 41599
rect 45097 41559 45155 41565
rect 45186 41556 45192 41608
rect 45244 41596 45250 41608
rect 48409 41599 48467 41605
rect 45244 41568 45289 41596
rect 45388 41568 47624 41596
rect 45244 41556 45250 41568
rect 39942 41528 39948 41540
rect 38488 41500 39948 41528
rect 21818 41460 21824 41472
rect 21192 41432 21824 41460
rect 21818 41420 21824 41432
rect 21876 41420 21882 41472
rect 23753 41463 23811 41469
rect 23753 41429 23765 41463
rect 23799 41460 23811 41463
rect 24578 41460 24584 41472
rect 23799 41432 24584 41460
rect 23799 41429 23811 41432
rect 23753 41423 23811 41429
rect 24578 41420 24584 41432
rect 24636 41420 24642 41472
rect 25038 41420 25044 41472
rect 25096 41460 25102 41472
rect 27157 41463 27215 41469
rect 27157 41460 27169 41463
rect 25096 41432 27169 41460
rect 25096 41420 25102 41432
rect 27157 41429 27169 41432
rect 27203 41429 27215 41463
rect 31938 41460 31944 41472
rect 31899 41432 31944 41460
rect 27157 41423 27215 41429
rect 31938 41420 31944 41432
rect 31996 41420 32002 41472
rect 32122 41420 32128 41472
rect 32180 41460 32186 41472
rect 32416 41460 32444 41491
rect 32600 41472 32628 41500
rect 39942 41488 39948 41500
rect 40000 41488 40006 41540
rect 42334 41488 42340 41540
rect 42392 41528 42398 41540
rect 42392 41500 42656 41528
rect 42392 41488 42398 41500
rect 42628 41472 42656 41500
rect 42886 41488 42892 41540
rect 42944 41528 42950 41540
rect 45388 41528 45416 41568
rect 42944 41500 45416 41528
rect 42944 41488 42950 41500
rect 47302 41488 47308 41540
rect 47360 41528 47366 41540
rect 47489 41531 47547 41537
rect 47489 41528 47501 41531
rect 47360 41500 47501 41528
rect 47360 41488 47366 41500
rect 47489 41497 47501 41500
rect 47535 41497 47547 41531
rect 47596 41528 47624 41568
rect 48409 41565 48421 41599
rect 48455 41596 48467 41599
rect 48498 41596 48504 41608
rect 48455 41568 48504 41596
rect 48455 41565 48467 41568
rect 48409 41559 48467 41565
rect 48498 41556 48504 41568
rect 48556 41596 48562 41608
rect 50062 41596 50068 41608
rect 48556 41568 50068 41596
rect 48556 41556 48562 41568
rect 50062 41556 50068 41568
rect 50120 41556 50126 41608
rect 50706 41596 50712 41608
rect 50667 41568 50712 41596
rect 50706 41556 50712 41568
rect 50764 41556 50770 41608
rect 51166 41596 51172 41608
rect 51127 41568 51172 41596
rect 51166 41556 51172 41568
rect 51224 41556 51230 41608
rect 51353 41599 51411 41605
rect 51353 41565 51365 41599
rect 51399 41596 51411 41599
rect 56965 41599 57023 41605
rect 51399 41568 51433 41596
rect 51399 41565 51411 41568
rect 51353 41559 51411 41565
rect 56965 41565 56977 41599
rect 57011 41596 57023 41599
rect 57238 41596 57244 41608
rect 57011 41568 57244 41596
rect 57011 41565 57023 41568
rect 56965 41559 57023 41565
rect 51368 41528 51396 41559
rect 57238 41556 57244 41568
rect 57296 41556 57302 41608
rect 52546 41528 52552 41540
rect 47596 41500 52552 41528
rect 47489 41491 47547 41497
rect 52546 41488 52552 41500
rect 52604 41488 52610 41540
rect 56689 41531 56747 41537
rect 56689 41497 56701 41531
rect 56735 41528 56747 41531
rect 57146 41528 57152 41540
rect 56735 41500 57152 41528
rect 56735 41497 56747 41500
rect 56689 41491 56747 41497
rect 57146 41488 57152 41500
rect 57204 41488 57210 41540
rect 32180 41432 32444 41460
rect 32180 41420 32186 41432
rect 32582 41420 32588 41472
rect 32640 41420 32646 41472
rect 33042 41420 33048 41472
rect 33100 41460 33106 41472
rect 33413 41463 33471 41469
rect 33413 41460 33425 41463
rect 33100 41432 33425 41460
rect 33100 41420 33106 41432
rect 33413 41429 33425 41432
rect 33459 41429 33471 41463
rect 33413 41423 33471 41429
rect 37461 41463 37519 41469
rect 37461 41429 37473 41463
rect 37507 41460 37519 41463
rect 38654 41460 38660 41472
rect 37507 41432 38660 41460
rect 37507 41429 37519 41432
rect 37461 41423 37519 41429
rect 38654 41420 38660 41432
rect 38712 41420 38718 41472
rect 42610 41420 42616 41472
rect 42668 41420 42674 41472
rect 45278 41460 45284 41472
rect 45239 41432 45284 41460
rect 45278 41420 45284 41432
rect 45336 41420 45342 41472
rect 47394 41420 47400 41472
rect 47452 41460 47458 41472
rect 47949 41463 48007 41469
rect 47949 41460 47961 41463
rect 47452 41432 47961 41460
rect 47452 41420 47458 41432
rect 47949 41429 47961 41432
rect 47995 41429 48007 41463
rect 47949 41423 48007 41429
rect 50525 41463 50583 41469
rect 50525 41429 50537 41463
rect 50571 41460 50583 41463
rect 50982 41460 50988 41472
rect 50571 41432 50988 41460
rect 50571 41429 50583 41432
rect 50525 41423 50583 41429
rect 50982 41420 50988 41432
rect 51040 41420 51046 41472
rect 51074 41420 51080 41472
rect 51132 41460 51138 41472
rect 51353 41463 51411 41469
rect 51353 41460 51365 41463
rect 51132 41432 51365 41460
rect 51132 41420 51138 41432
rect 51353 41429 51365 41432
rect 51399 41460 51411 41463
rect 51442 41460 51448 41472
rect 51399 41432 51448 41460
rect 51399 41429 51411 41432
rect 51353 41423 51411 41429
rect 51442 41420 51448 41432
rect 51500 41420 51506 41472
rect 56778 41420 56784 41472
rect 56836 41460 56842 41472
rect 56873 41463 56931 41469
rect 56873 41460 56885 41463
rect 56836 41432 56885 41460
rect 56836 41420 56842 41432
rect 56873 41429 56885 41432
rect 56919 41429 56931 41463
rect 56873 41423 56931 41429
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 22186 41256 22192 41268
rect 22147 41228 22192 41256
rect 22186 41216 22192 41228
rect 22244 41216 22250 41268
rect 24121 41259 24179 41265
rect 24121 41225 24133 41259
rect 24167 41256 24179 41259
rect 24854 41256 24860 41268
rect 24167 41228 24860 41256
rect 24167 41225 24179 41228
rect 24121 41219 24179 41225
rect 24854 41216 24860 41228
rect 24912 41216 24918 41268
rect 27522 41216 27528 41268
rect 27580 41256 27586 41268
rect 30834 41256 30840 41268
rect 27580 41228 30840 41256
rect 27580 41216 27586 41228
rect 30834 41216 30840 41228
rect 30892 41216 30898 41268
rect 33502 41256 33508 41268
rect 33463 41228 33508 41256
rect 33502 41216 33508 41228
rect 33560 41216 33566 41268
rect 33594 41216 33600 41268
rect 33652 41256 33658 41268
rect 34057 41259 34115 41265
rect 34057 41256 34069 41259
rect 33652 41228 34069 41256
rect 33652 41216 33658 41228
rect 34057 41225 34069 41228
rect 34103 41225 34115 41259
rect 34057 41219 34115 41225
rect 38194 41216 38200 41268
rect 38252 41256 38258 41268
rect 38289 41259 38347 41265
rect 38289 41256 38301 41259
rect 38252 41228 38301 41256
rect 38252 41216 38258 41228
rect 38289 41225 38301 41228
rect 38335 41225 38347 41259
rect 38289 41219 38347 41225
rect 39114 41216 39120 41268
rect 39172 41256 39178 41268
rect 39209 41259 39267 41265
rect 39209 41256 39221 41259
rect 39172 41228 39221 41256
rect 39172 41216 39178 41228
rect 39209 41225 39221 41228
rect 39255 41256 39267 41259
rect 39255 41228 39712 41256
rect 39255 41225 39267 41228
rect 39209 41219 39267 41225
rect 22738 41188 22744 41200
rect 20640 41160 22744 41188
rect 20640 41129 20668 41160
rect 22738 41148 22744 41160
rect 22796 41148 22802 41200
rect 29270 41148 29276 41200
rect 29328 41188 29334 41200
rect 32306 41188 32312 41200
rect 29328 41160 31754 41188
rect 32267 41160 32312 41188
rect 29328 41148 29334 41160
rect 20625 41123 20683 41129
rect 20625 41089 20637 41123
rect 20671 41089 20683 41123
rect 22005 41123 22063 41129
rect 22005 41120 22017 41123
rect 20625 41083 20683 41089
rect 21008 41092 22017 41120
rect 21008 41064 21036 41092
rect 22005 41089 22017 41092
rect 22051 41089 22063 41123
rect 23934 41120 23940 41132
rect 23895 41092 23940 41120
rect 22005 41083 22063 41089
rect 23934 41080 23940 41092
rect 23992 41080 23998 41132
rect 24118 41120 24124 41132
rect 24079 41092 24124 41120
rect 24118 41080 24124 41092
rect 24176 41080 24182 41132
rect 24578 41120 24584 41132
rect 24539 41092 24584 41120
rect 24578 41080 24584 41092
rect 24636 41080 24642 41132
rect 27893 41123 27951 41129
rect 27893 41089 27905 41123
rect 27939 41120 27951 41123
rect 29546 41120 29552 41132
rect 27939 41092 29552 41120
rect 27939 41089 27951 41092
rect 27893 41083 27951 41089
rect 29546 41080 29552 41092
rect 29604 41080 29610 41132
rect 29641 41123 29699 41129
rect 29641 41089 29653 41123
rect 29687 41089 29699 41123
rect 29822 41120 29828 41132
rect 29783 41092 29828 41120
rect 29641 41083 29699 41089
rect 20530 41052 20536 41064
rect 20491 41024 20536 41052
rect 20530 41012 20536 41024
rect 20588 41012 20594 41064
rect 20990 41052 20996 41064
rect 20951 41024 20996 41052
rect 20990 41012 20996 41024
rect 21048 41012 21054 41064
rect 21821 41055 21879 41061
rect 21821 41021 21833 41055
rect 21867 41052 21879 41055
rect 23658 41052 23664 41064
rect 21867 41024 23664 41052
rect 21867 41021 21879 41024
rect 21821 41015 21879 41021
rect 19978 40944 19984 40996
rect 20036 40984 20042 40996
rect 21836 40984 21864 41015
rect 23658 41012 23664 41024
rect 23716 41012 23722 41064
rect 24857 41055 24915 41061
rect 24857 41021 24869 41055
rect 24903 41052 24915 41055
rect 24946 41052 24952 41064
rect 24903 41024 24952 41052
rect 24903 41021 24915 41024
rect 24857 41015 24915 41021
rect 24946 41012 24952 41024
rect 25004 41052 25010 41064
rect 26418 41052 26424 41064
rect 25004 41024 26424 41052
rect 25004 41012 25010 41024
rect 26418 41012 26424 41024
rect 26476 41012 26482 41064
rect 27614 41052 27620 41064
rect 27575 41024 27620 41052
rect 27614 41012 27620 41024
rect 27672 41012 27678 41064
rect 29656 41052 29684 41083
rect 29822 41080 29828 41092
rect 29880 41080 29886 41132
rect 30190 41080 30196 41132
rect 30248 41120 30254 41132
rect 30285 41123 30343 41129
rect 30285 41120 30297 41123
rect 30248 41092 30297 41120
rect 30248 41080 30254 41092
rect 30285 41089 30297 41092
rect 30331 41089 30343 41123
rect 30285 41083 30343 41089
rect 30466 41080 30472 41132
rect 30524 41120 30530 41132
rect 30561 41123 30619 41129
rect 30561 41120 30573 41123
rect 30524 41092 30573 41120
rect 30524 41080 30530 41092
rect 30561 41089 30573 41092
rect 30607 41089 30619 41123
rect 30561 41083 30619 41089
rect 31386 41052 31392 41064
rect 29656 41024 31392 41052
rect 30208 40996 30236 41024
rect 31386 41012 31392 41024
rect 31444 41012 31450 41064
rect 24762 40984 24768 40996
rect 20036 40956 21864 40984
rect 24723 40956 24768 40984
rect 20036 40944 20042 40956
rect 24762 40944 24768 40956
rect 24820 40944 24826 40996
rect 29178 40944 29184 40996
rect 29236 40984 29242 40996
rect 30006 40984 30012 40996
rect 29236 40956 30012 40984
rect 29236 40944 29242 40956
rect 30006 40944 30012 40956
rect 30064 40944 30070 40996
rect 30190 40944 30196 40996
rect 30248 40944 30254 40996
rect 24670 40916 24676 40928
rect 24631 40888 24676 40916
rect 24670 40876 24676 40888
rect 24728 40876 24734 40928
rect 28350 40876 28356 40928
rect 28408 40916 28414 40928
rect 28629 40919 28687 40925
rect 28629 40916 28641 40919
rect 28408 40888 28641 40916
rect 28408 40876 28414 40888
rect 28629 40885 28641 40888
rect 28675 40885 28687 40919
rect 28629 40879 28687 40885
rect 29641 40919 29699 40925
rect 29641 40885 29653 40919
rect 29687 40916 29699 40919
rect 30742 40916 30748 40928
rect 29687 40888 30748 40916
rect 29687 40885 29699 40888
rect 29641 40879 29699 40885
rect 30742 40876 30748 40888
rect 30800 40876 30806 40928
rect 31726 40916 31754 41160
rect 32306 41148 32312 41160
rect 32364 41148 32370 41200
rect 32401 41191 32459 41197
rect 32401 41157 32413 41191
rect 32447 41188 32459 41191
rect 35618 41188 35624 41200
rect 32447 41160 35624 41188
rect 32447 41157 32459 41160
rect 32401 41151 32459 41157
rect 35618 41148 35624 41160
rect 35676 41148 35682 41200
rect 39684 41197 39712 41228
rect 39942 41216 39948 41268
rect 40000 41256 40006 41268
rect 40037 41259 40095 41265
rect 40037 41256 40049 41259
rect 40000 41228 40049 41256
rect 40000 41216 40006 41228
rect 40037 41225 40049 41228
rect 40083 41225 40095 41259
rect 40037 41219 40095 41225
rect 41601 41259 41659 41265
rect 41601 41225 41613 41259
rect 41647 41256 41659 41259
rect 41690 41256 41696 41268
rect 41647 41228 41696 41256
rect 41647 41225 41659 41228
rect 41601 41219 41659 41225
rect 41690 41216 41696 41228
rect 41748 41216 41754 41268
rect 43165 41259 43223 41265
rect 43165 41225 43177 41259
rect 43211 41256 43223 41259
rect 43438 41256 43444 41268
rect 43211 41228 43444 41256
rect 43211 41225 43223 41228
rect 43165 41219 43223 41225
rect 43438 41216 43444 41228
rect 43496 41216 43502 41268
rect 49234 41256 49240 41268
rect 46860 41228 49096 41256
rect 49195 41228 49240 41256
rect 39669 41191 39727 41197
rect 39669 41157 39681 41191
rect 39715 41157 39727 41191
rect 39669 41151 39727 41157
rect 39776 41160 41644 41188
rect 32122 41120 32128 41132
rect 32083 41092 32128 41120
rect 32122 41080 32128 41092
rect 32180 41080 32186 41132
rect 32493 41123 32551 41129
rect 32493 41089 32505 41123
rect 32539 41120 32551 41123
rect 32582 41120 32588 41132
rect 32539 41092 32588 41120
rect 32539 41089 32551 41092
rect 32493 41083 32551 41089
rect 32582 41080 32588 41092
rect 32640 41080 32646 41132
rect 33134 41120 33140 41132
rect 33095 41092 33140 41120
rect 33134 41080 33140 41092
rect 33192 41080 33198 41132
rect 33321 41123 33379 41129
rect 33321 41089 33333 41123
rect 33367 41120 33379 41123
rect 33410 41120 33416 41132
rect 33367 41092 33416 41120
rect 33367 41089 33379 41092
rect 33321 41083 33379 41089
rect 33410 41080 33416 41092
rect 33468 41080 33474 41132
rect 33965 41123 34023 41129
rect 33965 41089 33977 41123
rect 34011 41089 34023 41123
rect 34146 41120 34152 41132
rect 34107 41092 34152 41120
rect 33965 41083 34023 41089
rect 33980 41052 34008 41083
rect 34146 41080 34152 41092
rect 34204 41080 34210 41132
rect 37918 41080 37924 41132
rect 37976 41120 37982 41132
rect 38013 41123 38071 41129
rect 38013 41120 38025 41123
rect 37976 41092 38025 41120
rect 37976 41080 37982 41092
rect 38013 41089 38025 41092
rect 38059 41089 38071 41123
rect 38013 41083 38071 41089
rect 38289 41123 38347 41129
rect 38289 41089 38301 41123
rect 38335 41120 38347 41123
rect 38470 41120 38476 41132
rect 38335 41092 38476 41120
rect 38335 41089 38347 41092
rect 38289 41083 38347 41089
rect 38470 41080 38476 41092
rect 38528 41120 38534 41132
rect 39025 41123 39083 41129
rect 38528 41092 38976 41120
rect 38528 41080 38534 41092
rect 33980 41024 34014 41052
rect 31846 40944 31852 40996
rect 31904 40984 31910 40996
rect 33986 40984 34014 41024
rect 37826 41012 37832 41064
rect 37884 41052 37890 41064
rect 38841 41055 38899 41061
rect 38841 41052 38853 41055
rect 37884 41024 38853 41052
rect 37884 41012 37890 41024
rect 38841 41021 38853 41024
rect 38887 41021 38899 41055
rect 38948 41052 38976 41092
rect 39025 41089 39037 41123
rect 39071 41120 39083 41123
rect 39776 41120 39804 41160
rect 41616 41132 41644 41160
rect 39071 41092 39804 41120
rect 39853 41123 39911 41129
rect 39071 41089 39083 41092
rect 39025 41083 39083 41089
rect 39853 41089 39865 41123
rect 39899 41089 39911 41123
rect 39853 41083 39911 41089
rect 40589 41123 40647 41129
rect 40589 41089 40601 41123
rect 40635 41120 40647 41123
rect 40678 41120 40684 41132
rect 40635 41092 40684 41120
rect 40635 41089 40647 41092
rect 40589 41083 40647 41089
rect 39868 41052 39896 41083
rect 40678 41080 40684 41092
rect 40736 41080 40742 41132
rect 40773 41123 40831 41129
rect 40773 41089 40785 41123
rect 40819 41120 40831 41123
rect 41414 41120 41420 41132
rect 40819 41092 41420 41120
rect 40819 41089 40831 41092
rect 40773 41083 40831 41089
rect 41414 41080 41420 41092
rect 41472 41080 41478 41132
rect 41509 41123 41567 41129
rect 41509 41089 41521 41123
rect 41555 41089 41567 41123
rect 41509 41083 41567 41089
rect 38948 41024 39896 41052
rect 38841 41015 38899 41021
rect 31904 40956 34014 40984
rect 38856 40984 38884 41015
rect 40862 41012 40868 41064
rect 40920 41052 40926 41064
rect 41524 41052 41552 41083
rect 41598 41080 41604 41132
rect 41656 41080 41662 41132
rect 41693 41123 41751 41129
rect 41693 41089 41705 41123
rect 41739 41120 41751 41123
rect 41782 41120 41788 41132
rect 41739 41092 41788 41120
rect 41739 41089 41751 41092
rect 41693 41083 41751 41089
rect 41782 41080 41788 41092
rect 41840 41080 41846 41132
rect 42886 41120 42892 41132
rect 42847 41092 42892 41120
rect 42886 41080 42892 41092
rect 42944 41080 42950 41132
rect 42981 41123 43039 41129
rect 42981 41089 42993 41123
rect 43027 41089 43039 41123
rect 42981 41083 43039 41089
rect 40920 41024 41552 41052
rect 40920 41012 40926 41024
rect 42426 41012 42432 41064
rect 42484 41052 42490 41064
rect 42996 41052 43024 41083
rect 45922 41080 45928 41132
rect 45980 41120 45986 41132
rect 46290 41120 46296 41132
rect 45980 41092 46296 41120
rect 45980 41080 45986 41092
rect 46290 41080 46296 41092
rect 46348 41120 46354 41132
rect 46860 41129 46888 41228
rect 47118 41148 47124 41200
rect 47176 41188 47182 41200
rect 48041 41191 48099 41197
rect 48041 41188 48053 41191
rect 47176 41160 48053 41188
rect 47176 41148 47182 41160
rect 48041 41157 48053 41160
rect 48087 41188 48099 41191
rect 48869 41191 48927 41197
rect 48869 41188 48881 41191
rect 48087 41160 48881 41188
rect 48087 41157 48099 41160
rect 48041 41151 48099 41157
rect 48869 41157 48881 41160
rect 48915 41157 48927 41191
rect 49068 41188 49096 41228
rect 49234 41216 49240 41228
rect 49292 41216 49298 41268
rect 49881 41259 49939 41265
rect 49881 41225 49893 41259
rect 49927 41225 49939 41259
rect 49881 41219 49939 41225
rect 50065 41259 50123 41265
rect 50065 41225 50077 41259
rect 50111 41256 50123 41259
rect 51166 41256 51172 41268
rect 50111 41228 51172 41256
rect 50111 41225 50123 41228
rect 50065 41219 50123 41225
rect 49602 41188 49608 41200
rect 49068 41160 49608 41188
rect 48869 41151 48927 41157
rect 49602 41148 49608 41160
rect 49660 41148 49666 41200
rect 49896 41188 49924 41219
rect 51166 41216 51172 41228
rect 51224 41256 51230 41268
rect 51261 41259 51319 41265
rect 51261 41256 51273 41259
rect 51224 41228 51273 41256
rect 51224 41216 51230 41228
rect 51261 41225 51273 41228
rect 51307 41225 51319 41259
rect 51534 41256 51540 41268
rect 51495 41228 51540 41256
rect 51261 41219 51319 41225
rect 51534 41216 51540 41228
rect 51592 41216 51598 41268
rect 55306 41216 55312 41268
rect 55364 41256 55370 41268
rect 56321 41259 56379 41265
rect 56321 41256 56333 41259
rect 55364 41228 56333 41256
rect 55364 41216 55370 41228
rect 56321 41225 56333 41228
rect 56367 41225 56379 41259
rect 56321 41219 56379 41225
rect 57241 41259 57299 41265
rect 57241 41225 57253 41259
rect 57287 41256 57299 41259
rect 57330 41256 57336 41268
rect 57287 41228 57336 41256
rect 57287 41225 57299 41228
rect 57241 41219 57299 41225
rect 57330 41216 57336 41228
rect 57388 41216 57394 41268
rect 51902 41188 51908 41200
rect 49896 41160 51908 41188
rect 51902 41148 51908 41160
rect 51960 41148 51966 41200
rect 56778 41148 56784 41200
rect 56836 41188 56842 41200
rect 57146 41197 57152 41200
rect 56873 41191 56931 41197
rect 56873 41188 56885 41191
rect 56836 41160 56885 41188
rect 56836 41148 56842 41160
rect 56873 41157 56885 41160
rect 56919 41157 56931 41191
rect 56873 41151 56931 41157
rect 57089 41191 57152 41197
rect 57089 41157 57101 41191
rect 57135 41157 57152 41191
rect 57089 41151 57152 41157
rect 57146 41148 57152 41151
rect 57204 41148 57210 41200
rect 46845 41123 46903 41129
rect 46845 41120 46857 41123
rect 46348 41092 46857 41120
rect 46348 41080 46354 41092
rect 46845 41089 46857 41092
rect 46891 41089 46903 41123
rect 46845 41083 46903 41089
rect 47394 41080 47400 41132
rect 47452 41120 47458 41132
rect 47765 41123 47823 41129
rect 47765 41120 47777 41123
rect 47452 41092 47777 41120
rect 47452 41080 47458 41092
rect 47765 41089 47777 41092
rect 47811 41089 47823 41123
rect 47765 41083 47823 41089
rect 47858 41123 47916 41129
rect 47858 41089 47870 41123
rect 47904 41089 47916 41123
rect 47858 41083 47916 41089
rect 48133 41123 48191 41129
rect 48133 41089 48145 41123
rect 48179 41089 48191 41123
rect 48133 41083 48191 41089
rect 42484 41024 43024 41052
rect 42484 41012 42490 41024
rect 41690 40984 41696 40996
rect 38856 40956 41696 40984
rect 31904 40944 31910 40956
rect 41690 40944 41696 40956
rect 41748 40944 41754 40996
rect 42996 40984 43024 41024
rect 47210 41012 47216 41064
rect 47268 41052 47274 41064
rect 47872 41052 47900 41083
rect 47268 41024 47900 41052
rect 48148 41052 48176 41083
rect 48222 41080 48228 41132
rect 48280 41129 48286 41132
rect 48280 41120 48288 41129
rect 49053 41123 49111 41129
rect 48280 41092 48325 41120
rect 48280 41083 48288 41092
rect 49053 41089 49065 41123
rect 49099 41120 49111 41123
rect 49234 41120 49240 41132
rect 49099 41092 49240 41120
rect 49099 41089 49111 41092
rect 49053 41083 49111 41089
rect 48280 41080 48286 41083
rect 49234 41080 49240 41092
rect 49292 41080 49298 41132
rect 50062 41120 50068 41132
rect 49975 41092 50068 41120
rect 50062 41080 50068 41092
rect 50120 41120 50126 41132
rect 50982 41120 50988 41132
rect 50120 41092 50988 41120
rect 50120 41080 50126 41092
rect 50982 41080 50988 41092
rect 51040 41080 51046 41132
rect 51169 41123 51227 41129
rect 51169 41120 51181 41123
rect 51092 41092 51181 41120
rect 48682 41052 48688 41064
rect 48148 41024 48688 41052
rect 47268 41012 47274 41024
rect 48682 41012 48688 41024
rect 48740 41012 48746 41064
rect 49252 41052 49280 41080
rect 50522 41052 50528 41064
rect 49252 41024 50384 41052
rect 50483 41024 50528 41052
rect 49510 40984 49516 40996
rect 42996 40956 49516 40984
rect 49510 40944 49516 40956
rect 49568 40944 49574 40996
rect 50356 40984 50384 41024
rect 50522 41012 50528 41024
rect 50580 41012 50586 41064
rect 51092 40996 51120 41092
rect 51169 41089 51181 41092
rect 51215 41089 51227 41123
rect 51169 41083 51227 41089
rect 51353 41123 51411 41129
rect 51353 41089 51365 41123
rect 51399 41120 51411 41123
rect 51997 41123 52055 41129
rect 51399 41092 51856 41120
rect 51399 41089 51411 41092
rect 51353 41083 51411 41089
rect 51074 40984 51080 40996
rect 50356 40956 51080 40984
rect 51074 40944 51080 40956
rect 51132 40944 51138 40996
rect 51828 40984 51856 41092
rect 51997 41089 52009 41123
rect 52043 41089 52055 41123
rect 52178 41120 52184 41132
rect 52139 41092 52184 41120
rect 51997 41083 52055 41089
rect 52012 41052 52040 41083
rect 52178 41080 52184 41092
rect 52236 41080 52242 41132
rect 56226 41120 56232 41132
rect 56187 41092 56232 41120
rect 56226 41080 56232 41092
rect 56284 41080 56290 41132
rect 56413 41123 56471 41129
rect 56413 41089 56425 41123
rect 56459 41120 56471 41123
rect 57238 41120 57244 41132
rect 56459 41092 57244 41120
rect 56459 41089 56471 41092
rect 56413 41083 56471 41089
rect 57238 41080 57244 41092
rect 57296 41080 57302 41132
rect 52454 41052 52460 41064
rect 52012 41024 52460 41052
rect 52454 41012 52460 41024
rect 52512 41012 52518 41064
rect 52730 40984 52736 40996
rect 51828 40956 52736 40984
rect 52730 40944 52736 40956
rect 52788 40944 52794 40996
rect 32677 40919 32735 40925
rect 32677 40916 32689 40919
rect 31726 40888 32689 40916
rect 32677 40885 32689 40888
rect 32723 40885 32735 40919
rect 32677 40879 32735 40885
rect 38562 40876 38568 40928
rect 38620 40916 38626 40928
rect 40589 40919 40647 40925
rect 40589 40916 40601 40919
rect 38620 40888 40601 40916
rect 38620 40876 38626 40888
rect 40589 40885 40601 40888
rect 40635 40885 40647 40919
rect 46934 40916 46940 40928
rect 46895 40888 46940 40916
rect 40589 40879 40647 40885
rect 46934 40876 46940 40888
rect 46992 40876 46998 40928
rect 47394 40876 47400 40928
rect 47452 40916 47458 40928
rect 48409 40919 48467 40925
rect 48409 40916 48421 40919
rect 47452 40888 48421 40916
rect 47452 40876 47458 40888
rect 48409 40885 48421 40888
rect 48455 40885 48467 40919
rect 48409 40879 48467 40885
rect 49418 40876 49424 40928
rect 49476 40916 49482 40928
rect 50433 40919 50491 40925
rect 50433 40916 50445 40919
rect 49476 40888 50445 40916
rect 49476 40876 49482 40888
rect 50433 40885 50445 40888
rect 50479 40885 50491 40919
rect 50433 40879 50491 40885
rect 51626 40876 51632 40928
rect 51684 40916 51690 40928
rect 52089 40919 52147 40925
rect 52089 40916 52101 40919
rect 51684 40888 52101 40916
rect 51684 40876 51690 40888
rect 52089 40885 52101 40888
rect 52135 40885 52147 40919
rect 52089 40879 52147 40885
rect 57057 40919 57115 40925
rect 57057 40885 57069 40919
rect 57103 40916 57115 40919
rect 57238 40916 57244 40928
rect 57103 40888 57244 40916
rect 57103 40885 57115 40888
rect 57057 40879 57115 40885
rect 57238 40876 57244 40888
rect 57296 40876 57302 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 21082 40712 21088 40724
rect 21043 40684 21088 40712
rect 21082 40672 21088 40684
rect 21140 40672 21146 40724
rect 21177 40715 21235 40721
rect 21177 40681 21189 40715
rect 21223 40712 21235 40715
rect 21726 40712 21732 40724
rect 21223 40684 21732 40712
rect 21223 40681 21235 40684
rect 21177 40675 21235 40681
rect 21726 40672 21732 40684
rect 21784 40672 21790 40724
rect 21818 40672 21824 40724
rect 21876 40712 21882 40724
rect 29914 40712 29920 40724
rect 21876 40684 21921 40712
rect 29875 40684 29920 40712
rect 21876 40672 21882 40684
rect 29914 40672 29920 40684
rect 29972 40672 29978 40724
rect 31294 40712 31300 40724
rect 31255 40684 31300 40712
rect 31294 40672 31300 40684
rect 31352 40672 31358 40724
rect 31481 40715 31539 40721
rect 31481 40681 31493 40715
rect 31527 40712 31539 40715
rect 31754 40712 31760 40724
rect 31527 40684 31760 40712
rect 31527 40681 31539 40684
rect 31481 40675 31539 40681
rect 31754 40672 31760 40684
rect 31812 40672 31818 40724
rect 35069 40715 35127 40721
rect 35069 40712 35081 40715
rect 33336 40684 35081 40712
rect 21910 40644 21916 40656
rect 21284 40616 21916 40644
rect 21284 40585 21312 40616
rect 21910 40604 21916 40616
rect 21968 40604 21974 40656
rect 22646 40604 22652 40656
rect 22704 40644 22710 40656
rect 24397 40647 24455 40653
rect 24397 40644 24409 40647
rect 22704 40616 24409 40644
rect 22704 40604 22710 40616
rect 24397 40613 24409 40616
rect 24443 40613 24455 40647
rect 24397 40607 24455 40613
rect 31386 40604 31392 40656
rect 31444 40644 31450 40656
rect 33336 40644 33364 40684
rect 34900 40656 34928 40684
rect 35069 40681 35081 40684
rect 35115 40681 35127 40715
rect 35069 40675 35127 40681
rect 37001 40715 37059 40721
rect 37001 40681 37013 40715
rect 37047 40712 37059 40715
rect 37274 40712 37280 40724
rect 37047 40684 37280 40712
rect 37047 40681 37059 40684
rect 37001 40675 37059 40681
rect 37274 40672 37280 40684
rect 37332 40672 37338 40724
rect 40770 40672 40776 40724
rect 40828 40712 40834 40724
rect 42153 40715 42211 40721
rect 42153 40712 42165 40715
rect 40828 40684 42165 40712
rect 40828 40672 40834 40684
rect 42153 40681 42165 40684
rect 42199 40681 42211 40715
rect 42153 40675 42211 40681
rect 42702 40672 42708 40724
rect 42760 40712 42766 40724
rect 47213 40715 47271 40721
rect 47213 40712 47225 40715
rect 42760 40684 47225 40712
rect 42760 40672 42766 40684
rect 47213 40681 47225 40684
rect 47259 40681 47271 40715
rect 47213 40675 47271 40681
rect 47946 40672 47952 40724
rect 48004 40712 48010 40724
rect 48409 40715 48467 40721
rect 48409 40712 48421 40715
rect 48004 40684 48421 40712
rect 48004 40672 48010 40684
rect 48409 40681 48421 40684
rect 48455 40681 48467 40715
rect 49510 40712 49516 40724
rect 49471 40684 49516 40712
rect 48409 40675 48467 40681
rect 49510 40672 49516 40684
rect 49568 40672 49574 40724
rect 49602 40672 49608 40724
rect 49660 40712 49666 40724
rect 52454 40712 52460 40724
rect 49660 40684 52460 40712
rect 49660 40672 49666 40684
rect 52454 40672 52460 40684
rect 52512 40672 52518 40724
rect 56226 40672 56232 40724
rect 56284 40712 56290 40724
rect 56689 40715 56747 40721
rect 56689 40712 56701 40715
rect 56284 40684 56701 40712
rect 56284 40672 56290 40684
rect 56689 40681 56701 40684
rect 56735 40681 56747 40715
rect 57238 40712 57244 40724
rect 57199 40684 57244 40712
rect 56689 40675 56747 40681
rect 57238 40672 57244 40684
rect 57296 40672 57302 40724
rect 31444 40616 33364 40644
rect 33505 40647 33563 40653
rect 31444 40604 31450 40616
rect 33505 40613 33517 40647
rect 33551 40644 33563 40647
rect 33870 40644 33876 40656
rect 33551 40616 33876 40644
rect 33551 40613 33563 40616
rect 33505 40607 33563 40613
rect 33870 40604 33876 40616
rect 33928 40604 33934 40656
rect 34882 40604 34888 40656
rect 34940 40604 34946 40656
rect 39853 40647 39911 40653
rect 39853 40644 39865 40647
rect 38856 40616 39865 40644
rect 21269 40579 21327 40585
rect 21269 40545 21281 40579
rect 21315 40545 21327 40579
rect 22278 40576 22284 40588
rect 21269 40539 21327 40545
rect 21744 40548 22284 40576
rect 21744 40517 21772 40548
rect 22278 40536 22284 40548
rect 22336 40536 22342 40588
rect 23658 40536 23664 40588
rect 23716 40576 23722 40588
rect 24486 40576 24492 40588
rect 23716 40548 24492 40576
rect 23716 40536 23722 40548
rect 24486 40536 24492 40548
rect 24544 40576 24550 40588
rect 24765 40579 24823 40585
rect 24765 40576 24777 40579
rect 24544 40548 24777 40576
rect 24544 40536 24550 40548
rect 24765 40545 24777 40548
rect 24811 40545 24823 40579
rect 24765 40539 24823 40545
rect 27982 40536 27988 40588
rect 28040 40576 28046 40588
rect 28169 40579 28227 40585
rect 28169 40576 28181 40579
rect 28040 40548 28181 40576
rect 28040 40536 28046 40548
rect 28169 40545 28181 40548
rect 28215 40545 28227 40579
rect 28169 40539 28227 40545
rect 30098 40536 30104 40588
rect 30156 40576 30162 40588
rect 30469 40579 30527 40585
rect 30469 40576 30481 40579
rect 30156 40548 30481 40576
rect 30156 40536 30162 40548
rect 30469 40545 30481 40548
rect 30515 40545 30527 40579
rect 31754 40576 31760 40588
rect 30469 40539 30527 40545
rect 31588 40548 31760 40576
rect 20993 40511 21051 40517
rect 20993 40477 21005 40511
rect 21039 40477 21051 40511
rect 20993 40471 21051 40477
rect 21729 40511 21787 40517
rect 21729 40477 21741 40511
rect 21775 40477 21787 40511
rect 21910 40508 21916 40520
rect 21871 40480 21916 40508
rect 21729 40471 21787 40477
rect 21008 40440 21036 40471
rect 21910 40468 21916 40480
rect 21968 40468 21974 40520
rect 24302 40468 24308 40520
rect 24360 40508 24366 40520
rect 24581 40511 24639 40517
rect 24581 40508 24593 40511
rect 24360 40480 24593 40508
rect 24360 40468 24366 40480
rect 24581 40477 24593 40480
rect 24627 40477 24639 40511
rect 24581 40471 24639 40477
rect 24857 40511 24915 40517
rect 24857 40477 24869 40511
rect 24903 40508 24915 40511
rect 25406 40508 25412 40520
rect 24903 40480 25412 40508
rect 24903 40477 24915 40480
rect 24857 40471 24915 40477
rect 25406 40468 25412 40480
rect 25464 40468 25470 40520
rect 27709 40511 27767 40517
rect 27709 40477 27721 40511
rect 27755 40477 27767 40511
rect 28350 40508 28356 40520
rect 28311 40480 28356 40508
rect 27709 40471 27767 40477
rect 22186 40440 22192 40452
rect 21008 40412 22192 40440
rect 22186 40400 22192 40412
rect 22244 40400 22250 40452
rect 22738 40400 22744 40452
rect 22796 40440 22802 40452
rect 23201 40443 23259 40449
rect 23201 40440 23213 40443
rect 22796 40412 23213 40440
rect 22796 40400 22802 40412
rect 23201 40409 23213 40412
rect 23247 40440 23259 40443
rect 23750 40440 23756 40452
rect 23247 40412 23756 40440
rect 23247 40409 23259 40412
rect 23201 40403 23259 40409
rect 23750 40400 23756 40412
rect 23808 40440 23814 40452
rect 25317 40443 25375 40449
rect 25317 40440 25329 40443
rect 23808 40412 25329 40440
rect 23808 40400 23814 40412
rect 25317 40409 25329 40412
rect 25363 40409 25375 40443
rect 25498 40440 25504 40452
rect 25459 40412 25504 40440
rect 25317 40403 25375 40409
rect 25498 40400 25504 40412
rect 25556 40400 25562 40452
rect 27724 40440 27752 40471
rect 28350 40468 28356 40480
rect 28408 40468 28414 40520
rect 30377 40511 30435 40517
rect 30377 40477 30389 40511
rect 30423 40508 30435 40511
rect 31588 40508 31616 40548
rect 31754 40536 31760 40548
rect 31812 40536 31818 40588
rect 31941 40579 31999 40585
rect 31941 40545 31953 40579
rect 31987 40576 31999 40579
rect 33134 40576 33140 40588
rect 31987 40548 33140 40576
rect 31987 40545 31999 40548
rect 31941 40539 31999 40545
rect 30423 40480 31616 40508
rect 30423 40477 30435 40480
rect 30377 40471 30435 40477
rect 31662 40468 31668 40520
rect 31720 40508 31726 40520
rect 31956 40508 31984 40539
rect 33134 40536 33140 40548
rect 33192 40536 33198 40588
rect 37826 40576 37832 40588
rect 34900 40548 37832 40576
rect 31720 40480 31984 40508
rect 32217 40511 32275 40517
rect 31720 40468 31726 40480
rect 32217 40477 32229 40511
rect 32263 40508 32275 40511
rect 32490 40508 32496 40520
rect 32263 40480 32496 40508
rect 32263 40477 32275 40480
rect 32217 40471 32275 40477
rect 32490 40468 32496 40480
rect 32548 40468 32554 40520
rect 32674 40468 32680 40520
rect 32732 40508 32738 40520
rect 33321 40511 33379 40517
rect 33321 40508 33333 40511
rect 32732 40480 33333 40508
rect 32732 40468 32738 40480
rect 33321 40477 33333 40480
rect 33367 40508 33379 40511
rect 33594 40508 33600 40520
rect 33367 40480 33600 40508
rect 33367 40477 33379 40480
rect 33321 40471 33379 40477
rect 33594 40468 33600 40480
rect 33652 40468 33658 40520
rect 34900 40517 34928 40548
rect 37826 40536 37832 40548
rect 37884 40536 37890 40588
rect 37918 40536 37924 40588
rect 37976 40576 37982 40588
rect 38856 40585 38884 40616
rect 39853 40613 39865 40616
rect 39899 40613 39911 40647
rect 39853 40607 39911 40613
rect 40218 40604 40224 40656
rect 40276 40644 40282 40656
rect 40276 40616 46980 40644
rect 40276 40604 40282 40616
rect 38841 40579 38899 40585
rect 37976 40548 38792 40576
rect 37976 40536 37982 40548
rect 34885 40511 34943 40517
rect 34885 40477 34897 40511
rect 34931 40477 34943 40511
rect 34885 40471 34943 40477
rect 35161 40511 35219 40517
rect 35161 40477 35173 40511
rect 35207 40477 35219 40511
rect 35161 40471 35219 40477
rect 37001 40511 37059 40517
rect 37001 40477 37013 40511
rect 37047 40508 37059 40511
rect 37047 40480 37136 40508
rect 37047 40477 37059 40480
rect 37001 40471 37059 40477
rect 28537 40443 28595 40449
rect 28537 40440 28549 40443
rect 27724 40412 28549 40440
rect 28537 40409 28549 40412
rect 28583 40409 28595 40443
rect 31110 40440 31116 40452
rect 31071 40412 31116 40440
rect 28537 40403 28595 40409
rect 31110 40400 31116 40412
rect 31168 40400 31174 40452
rect 32582 40400 32588 40452
rect 32640 40440 32646 40452
rect 34974 40440 34980 40452
rect 32640 40412 34980 40440
rect 32640 40400 32646 40412
rect 34974 40400 34980 40412
rect 35032 40440 35038 40452
rect 35176 40440 35204 40471
rect 35032 40412 35204 40440
rect 37108 40440 37136 40480
rect 37182 40468 37188 40520
rect 37240 40508 37246 40520
rect 38562 40508 38568 40520
rect 37240 40480 37285 40508
rect 38523 40480 38568 40508
rect 37240 40468 37246 40480
rect 38562 40468 38568 40480
rect 38620 40468 38626 40520
rect 38764 40517 38792 40548
rect 38841 40545 38853 40579
rect 38887 40545 38899 40579
rect 38841 40539 38899 40545
rect 39942 40536 39948 40588
rect 40000 40576 40006 40588
rect 40037 40579 40095 40585
rect 40037 40576 40049 40579
rect 40000 40548 40049 40576
rect 40000 40536 40006 40548
rect 40037 40545 40049 40548
rect 40083 40545 40095 40579
rect 40037 40539 40095 40545
rect 40405 40579 40463 40585
rect 40405 40545 40417 40579
rect 40451 40576 40463 40579
rect 40862 40576 40868 40588
rect 40451 40548 40868 40576
rect 40451 40545 40463 40548
rect 40405 40539 40463 40545
rect 40862 40536 40868 40548
rect 40920 40536 40926 40588
rect 43073 40579 43131 40585
rect 43073 40576 43085 40579
rect 41800 40548 43085 40576
rect 38749 40511 38807 40517
rect 38749 40477 38761 40511
rect 38795 40477 38807 40511
rect 38749 40471 38807 40477
rect 38933 40511 38991 40517
rect 38933 40477 38945 40511
rect 38979 40477 38991 40511
rect 39114 40508 39120 40520
rect 39075 40480 39120 40508
rect 38933 40471 38991 40477
rect 38948 40440 38976 40471
rect 39114 40468 39120 40480
rect 39172 40508 39178 40520
rect 40129 40511 40187 40517
rect 39172 40480 40080 40508
rect 39172 40468 39178 40480
rect 40052 40440 40080 40480
rect 40129 40477 40141 40511
rect 40175 40508 40187 40511
rect 41049 40511 41107 40517
rect 41049 40508 41061 40511
rect 40175 40480 41061 40508
rect 40175 40477 40187 40480
rect 40129 40471 40187 40477
rect 41049 40477 41061 40480
rect 41095 40477 41107 40511
rect 41049 40471 41107 40477
rect 41233 40511 41291 40517
rect 41233 40477 41245 40511
rect 41279 40508 41291 40511
rect 41509 40511 41567 40517
rect 41279 40480 41414 40508
rect 41279 40477 41291 40480
rect 41233 40471 41291 40477
rect 40497 40443 40555 40449
rect 40497 40440 40509 40443
rect 37108 40412 39988 40440
rect 40052 40412 40509 40440
rect 35032 40400 35038 40412
rect 22278 40332 22284 40384
rect 22336 40372 22342 40384
rect 23293 40375 23351 40381
rect 23293 40372 23305 40375
rect 22336 40344 23305 40372
rect 22336 40332 22342 40344
rect 23293 40341 23305 40344
rect 23339 40341 23351 40375
rect 23293 40335 23351 40341
rect 25685 40375 25743 40381
rect 25685 40341 25697 40375
rect 25731 40372 25743 40375
rect 26234 40372 26240 40384
rect 25731 40344 26240 40372
rect 25731 40341 25743 40344
rect 25685 40335 25743 40341
rect 26234 40332 26240 40344
rect 26292 40332 26298 40384
rect 27525 40375 27583 40381
rect 27525 40341 27537 40375
rect 27571 40372 27583 40375
rect 27890 40372 27896 40384
rect 27571 40344 27896 40372
rect 27571 40341 27583 40344
rect 27525 40335 27583 40341
rect 27890 40332 27896 40344
rect 27948 40332 27954 40384
rect 30285 40375 30343 40381
rect 30285 40341 30297 40375
rect 30331 40372 30343 40375
rect 30374 40372 30380 40384
rect 30331 40344 30380 40372
rect 30331 40341 30343 40344
rect 30285 40335 30343 40341
rect 30374 40332 30380 40344
rect 30432 40332 30438 40384
rect 30466 40332 30472 40384
rect 30524 40372 30530 40384
rect 31313 40375 31371 40381
rect 31313 40372 31325 40375
rect 30524 40344 31325 40372
rect 30524 40332 30530 40344
rect 31313 40341 31325 40344
rect 31359 40341 31371 40375
rect 31313 40335 31371 40341
rect 33134 40332 33140 40384
rect 33192 40372 33198 40384
rect 33870 40372 33876 40384
rect 33192 40344 33876 40372
rect 33192 40332 33198 40344
rect 33870 40332 33876 40344
rect 33928 40332 33934 40384
rect 34701 40375 34759 40381
rect 34701 40341 34713 40375
rect 34747 40372 34759 40375
rect 34790 40372 34796 40384
rect 34747 40344 34796 40372
rect 34747 40341 34759 40344
rect 34701 40335 34759 40341
rect 34790 40332 34796 40344
rect 34848 40332 34854 40384
rect 37182 40332 37188 40384
rect 37240 40372 37246 40384
rect 38746 40372 38752 40384
rect 37240 40344 38752 40372
rect 37240 40332 37246 40344
rect 38746 40332 38752 40344
rect 38804 40372 38810 40384
rect 39114 40372 39120 40384
rect 38804 40344 39120 40372
rect 38804 40332 38810 40344
rect 39114 40332 39120 40344
rect 39172 40332 39178 40384
rect 39301 40375 39359 40381
rect 39301 40341 39313 40375
rect 39347 40372 39359 40375
rect 39482 40372 39488 40384
rect 39347 40344 39488 40372
rect 39347 40341 39359 40344
rect 39301 40335 39359 40341
rect 39482 40332 39488 40344
rect 39540 40332 39546 40384
rect 39960 40372 39988 40412
rect 40497 40409 40509 40412
rect 40543 40409 40555 40443
rect 41386 40440 41414 40480
rect 41509 40477 41521 40511
rect 41555 40508 41567 40511
rect 41598 40508 41604 40520
rect 41555 40480 41604 40508
rect 41555 40477 41567 40480
rect 41509 40471 41567 40477
rect 41598 40468 41604 40480
rect 41656 40468 41662 40520
rect 41690 40468 41696 40520
rect 41748 40517 41754 40520
rect 41748 40511 41763 40517
rect 41751 40508 41763 40511
rect 41800 40508 41828 40548
rect 43073 40545 43085 40548
rect 43119 40576 43131 40579
rect 43162 40576 43168 40588
rect 43119 40548 43168 40576
rect 43119 40545 43131 40548
rect 43073 40539 43131 40545
rect 43162 40536 43168 40548
rect 43220 40536 43226 40588
rect 46569 40579 46627 40585
rect 46569 40545 46581 40579
rect 46615 40576 46627 40579
rect 46842 40576 46848 40588
rect 46615 40548 46848 40576
rect 46615 40545 46627 40548
rect 46569 40539 46627 40545
rect 46842 40536 46848 40548
rect 46900 40536 46906 40588
rect 42150 40508 42156 40520
rect 41751 40480 41841 40508
rect 42111 40480 42156 40508
rect 41751 40477 41763 40480
rect 41748 40471 41763 40477
rect 41748 40468 41754 40471
rect 42150 40468 42156 40480
rect 42208 40468 42214 40520
rect 42242 40468 42248 40520
rect 42300 40508 42306 40520
rect 42337 40511 42395 40517
rect 42337 40508 42349 40511
rect 42300 40480 42349 40508
rect 42300 40468 42306 40480
rect 42337 40477 42349 40480
rect 42383 40477 42395 40511
rect 42886 40508 42892 40520
rect 42847 40480 42892 40508
rect 42337 40471 42395 40477
rect 42886 40468 42892 40480
rect 42944 40468 42950 40520
rect 46658 40468 46664 40520
rect 46716 40511 46722 40520
rect 46716 40505 46755 40511
rect 46743 40471 46755 40505
rect 46716 40468 46755 40471
rect 46697 40465 46755 40468
rect 42702 40440 42708 40452
rect 41386 40412 42708 40440
rect 40497 40403 40555 40409
rect 42702 40400 42708 40412
rect 42760 40400 42766 40452
rect 45186 40400 45192 40452
rect 45244 40440 45250 40452
rect 46293 40443 46351 40449
rect 46293 40440 46305 40443
rect 45244 40412 46305 40440
rect 45244 40400 45250 40412
rect 46293 40409 46305 40412
rect 46339 40409 46351 40443
rect 46474 40440 46480 40452
rect 46435 40412 46480 40440
rect 46293 40403 46351 40409
rect 46474 40400 46480 40412
rect 46532 40400 46538 40452
rect 46566 40400 46572 40452
rect 46624 40440 46630 40452
rect 46952 40440 46980 40616
rect 47578 40604 47584 40656
rect 47636 40644 47642 40656
rect 47854 40644 47860 40656
rect 47636 40616 47860 40644
rect 47636 40604 47642 40616
rect 47854 40604 47860 40616
rect 47912 40644 47918 40656
rect 47912 40616 49464 40644
rect 47912 40604 47918 40616
rect 48406 40576 48412 40588
rect 47596 40548 48412 40576
rect 47394 40508 47400 40520
rect 47355 40480 47400 40508
rect 47394 40468 47400 40480
rect 47452 40468 47458 40520
rect 47596 40517 47624 40548
rect 48406 40536 48412 40548
rect 48464 40536 48470 40588
rect 47581 40511 47639 40517
rect 47581 40477 47593 40511
rect 47627 40477 47639 40511
rect 47854 40508 47860 40520
rect 47815 40480 47860 40508
rect 47581 40471 47639 40477
rect 47854 40468 47860 40480
rect 47912 40468 47918 40520
rect 47946 40468 47952 40520
rect 48004 40508 48010 40520
rect 48317 40511 48375 40517
rect 48317 40508 48329 40511
rect 48004 40480 48329 40508
rect 48004 40468 48010 40480
rect 48317 40477 48329 40480
rect 48363 40477 48375 40511
rect 48317 40471 48375 40477
rect 48501 40511 48559 40517
rect 48501 40477 48513 40511
rect 48547 40508 48559 40511
rect 49326 40508 49332 40520
rect 48547 40480 49332 40508
rect 48547 40477 48559 40480
rect 48501 40471 48559 40477
rect 49326 40468 49332 40480
rect 49384 40468 49390 40520
rect 49436 40508 49464 40616
rect 49878 40604 49884 40656
rect 49936 40644 49942 40656
rect 50433 40647 50491 40653
rect 50433 40644 50445 40647
rect 49936 40616 50445 40644
rect 49936 40604 49942 40616
rect 50433 40613 50445 40616
rect 50479 40644 50491 40647
rect 51534 40644 51540 40656
rect 50479 40616 51540 40644
rect 50479 40613 50491 40616
rect 50433 40607 50491 40613
rect 51534 40604 51540 40616
rect 51592 40604 51598 40656
rect 50062 40536 50068 40588
rect 50120 40576 50126 40588
rect 50522 40576 50528 40588
rect 50120 40548 50528 40576
rect 50120 40536 50126 40548
rect 50356 40517 50384 40548
rect 50522 40536 50528 40548
rect 50580 40536 50586 40588
rect 51626 40576 51632 40588
rect 51587 40548 51632 40576
rect 51626 40536 51632 40548
rect 51684 40536 51690 40588
rect 50157 40511 50215 40517
rect 50157 40508 50169 40511
rect 49436 40480 50169 40508
rect 50157 40477 50169 40480
rect 50203 40477 50215 40511
rect 50157 40471 50215 40477
rect 50341 40511 50399 40517
rect 50341 40477 50353 40511
rect 50387 40477 50399 40511
rect 50341 40471 50399 40477
rect 51442 40468 51448 40520
rect 51500 40508 51506 40520
rect 51537 40511 51595 40517
rect 51537 40508 51549 40511
rect 51500 40480 51549 40508
rect 51500 40468 51506 40480
rect 51537 40477 51549 40480
rect 51583 40477 51595 40511
rect 51537 40471 51595 40477
rect 52365 40511 52423 40517
rect 52365 40477 52377 40511
rect 52411 40508 52423 40511
rect 52730 40508 52736 40520
rect 52411 40480 52736 40508
rect 52411 40477 52423 40480
rect 52365 40471 52423 40477
rect 52730 40468 52736 40480
rect 52788 40468 52794 40520
rect 55490 40508 55496 40520
rect 55451 40480 55496 40508
rect 55490 40468 55496 40480
rect 55548 40468 55554 40520
rect 55766 40508 55772 40520
rect 55727 40480 55772 40508
rect 55766 40468 55772 40480
rect 55824 40468 55830 40520
rect 56321 40511 56379 40517
rect 56321 40477 56333 40511
rect 56367 40508 56379 40511
rect 56410 40508 56416 40520
rect 56367 40480 56416 40508
rect 56367 40477 56379 40480
rect 56321 40471 56379 40477
rect 56410 40468 56416 40480
rect 56468 40508 56474 40520
rect 57149 40511 57207 40517
rect 57149 40508 57161 40511
rect 56468 40480 57161 40508
rect 56468 40468 56474 40480
rect 57149 40477 57161 40480
rect 57195 40477 57207 40511
rect 57149 40471 57207 40477
rect 57333 40511 57391 40517
rect 57333 40477 57345 40511
rect 57379 40477 57391 40511
rect 57333 40471 57391 40477
rect 47486 40440 47492 40452
rect 46624 40412 46669 40440
rect 46952 40412 47348 40440
rect 47447 40412 47492 40440
rect 46624 40400 46630 40412
rect 40402 40372 40408 40384
rect 39960 40344 40408 40372
rect 40402 40332 40408 40344
rect 40460 40332 40466 40384
rect 40586 40332 40592 40384
rect 40644 40372 40650 40384
rect 41506 40372 41512 40384
rect 40644 40344 41512 40372
rect 40644 40332 40650 40344
rect 41506 40332 41512 40344
rect 41564 40332 41570 40384
rect 47320 40372 47348 40412
rect 47486 40400 47492 40412
rect 47544 40400 47550 40452
rect 47670 40400 47676 40452
rect 47728 40449 47734 40452
rect 47728 40443 47757 40449
rect 47745 40440 47757 40443
rect 48130 40440 48136 40452
rect 47745 40412 48136 40440
rect 47745 40409 47757 40412
rect 47728 40403 47757 40409
rect 47728 40400 47734 40403
rect 48130 40400 48136 40412
rect 48188 40400 48194 40452
rect 49421 40443 49479 40449
rect 49421 40409 49433 40443
rect 49467 40440 49479 40443
rect 51166 40440 51172 40452
rect 49467 40412 51172 40440
rect 49467 40409 49479 40412
rect 49421 40403 49479 40409
rect 51166 40400 51172 40412
rect 51224 40400 51230 40452
rect 52178 40440 52184 40452
rect 51368 40412 52184 40440
rect 51258 40372 51264 40384
rect 47320 40344 51264 40372
rect 51258 40332 51264 40344
rect 51316 40372 51322 40384
rect 51368 40372 51396 40412
rect 52178 40400 52184 40412
rect 52236 40400 52242 40452
rect 54754 40400 54760 40452
rect 54812 40440 54818 40452
rect 55677 40443 55735 40449
rect 55677 40440 55689 40443
rect 54812 40412 55689 40440
rect 54812 40400 54818 40412
rect 55677 40409 55689 40412
rect 55723 40409 55735 40443
rect 55677 40403 55735 40409
rect 56226 40400 56232 40452
rect 56284 40440 56290 40452
rect 56505 40443 56563 40449
rect 56505 40440 56517 40443
rect 56284 40412 56517 40440
rect 56284 40400 56290 40412
rect 56505 40409 56517 40412
rect 56551 40440 56563 40443
rect 57348 40440 57376 40471
rect 56551 40412 57376 40440
rect 56551 40409 56563 40412
rect 56505 40403 56563 40409
rect 51902 40372 51908 40384
rect 51316 40344 51396 40372
rect 51863 40344 51908 40372
rect 51316 40332 51322 40344
rect 51902 40332 51908 40344
rect 51960 40332 51966 40384
rect 52454 40332 52460 40384
rect 52512 40372 52518 40384
rect 52549 40375 52607 40381
rect 52549 40372 52561 40375
rect 52512 40344 52561 40372
rect 52512 40332 52518 40344
rect 52549 40341 52561 40344
rect 52595 40341 52607 40375
rect 55306 40372 55312 40384
rect 55267 40344 55312 40372
rect 52549 40335 52607 40341
rect 55306 40332 55312 40344
rect 55364 40332 55370 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 23934 40168 23940 40180
rect 23895 40140 23940 40168
rect 23934 40128 23940 40140
rect 23992 40128 23998 40180
rect 25406 40168 25412 40180
rect 24044 40140 25412 40168
rect 20530 40060 20536 40112
rect 20588 40100 20594 40112
rect 22278 40100 22284 40112
rect 20588 40072 22284 40100
rect 20588 40060 20594 40072
rect 22278 40060 22284 40072
rect 22336 40060 22342 40112
rect 24044 40100 24072 40140
rect 25406 40128 25412 40140
rect 25464 40128 25470 40180
rect 25498 40128 25504 40180
rect 25556 40168 25562 40180
rect 25777 40171 25835 40177
rect 25777 40168 25789 40171
rect 25556 40140 25789 40168
rect 25556 40128 25562 40140
rect 25777 40137 25789 40140
rect 25823 40137 25835 40171
rect 25777 40131 25835 40137
rect 30101 40171 30159 40177
rect 30101 40137 30113 40171
rect 30147 40168 30159 40171
rect 30190 40168 30196 40180
rect 30147 40140 30196 40168
rect 30147 40137 30159 40140
rect 30101 40131 30159 40137
rect 30190 40128 30196 40140
rect 30248 40128 30254 40180
rect 30374 40128 30380 40180
rect 30432 40168 30438 40180
rect 31662 40168 31668 40180
rect 30432 40140 31668 40168
rect 30432 40128 30438 40140
rect 31662 40128 31668 40140
rect 31720 40168 31726 40180
rect 37918 40168 37924 40180
rect 31720 40128 31754 40168
rect 37879 40140 37924 40168
rect 37918 40128 37924 40140
rect 37976 40128 37982 40180
rect 38470 40168 38476 40180
rect 38431 40140 38476 40168
rect 38470 40128 38476 40140
rect 38528 40128 38534 40180
rect 40678 40128 40684 40180
rect 40736 40168 40742 40180
rect 40957 40171 41015 40177
rect 40957 40168 40969 40171
rect 40736 40140 40969 40168
rect 40736 40128 40742 40140
rect 40957 40137 40969 40140
rect 41003 40137 41015 40171
rect 40957 40131 41015 40137
rect 46934 40128 46940 40180
rect 46992 40168 46998 40180
rect 47670 40168 47676 40180
rect 46992 40140 47676 40168
rect 46992 40128 46998 40140
rect 47670 40128 47676 40140
rect 47728 40128 47734 40180
rect 48866 40168 48872 40180
rect 48056 40140 48872 40168
rect 23584 40072 24072 40100
rect 22186 39992 22192 40044
rect 22244 40032 22250 40044
rect 22465 40035 22523 40041
rect 22465 40032 22477 40035
rect 22244 40004 22477 40032
rect 22244 39992 22250 40004
rect 22465 40001 22477 40004
rect 22511 40032 22523 40035
rect 22830 40032 22836 40044
rect 22511 40004 22836 40032
rect 22511 40001 22523 40004
rect 22465 39995 22523 40001
rect 22830 39992 22836 40004
rect 22888 39992 22894 40044
rect 23584 40041 23612 40072
rect 24302 40060 24308 40112
rect 24360 40100 24366 40112
rect 29362 40100 29368 40112
rect 24360 40072 26464 40100
rect 24360 40060 24366 40072
rect 23569 40035 23627 40041
rect 23569 40001 23581 40035
rect 23615 40001 23627 40035
rect 23569 39995 23627 40001
rect 24486 39992 24492 40044
rect 24544 40032 24550 40044
rect 24653 40035 24711 40041
rect 24653 40032 24665 40035
rect 24544 40004 24665 40032
rect 24544 39992 24550 40004
rect 24653 40001 24665 40004
rect 24699 40001 24711 40035
rect 26234 40032 26240 40044
rect 26195 40004 26240 40032
rect 24653 39995 24711 40001
rect 26234 39992 26240 40004
rect 26292 39992 26298 40044
rect 26436 40041 26464 40072
rect 28184 40072 29368 40100
rect 26421 40035 26479 40041
rect 26421 40001 26433 40035
rect 26467 40001 26479 40035
rect 26421 39995 26479 40001
rect 27614 39992 27620 40044
rect 27672 40032 27678 40044
rect 28184 40041 28212 40072
rect 29362 40060 29368 40072
rect 29420 40060 29426 40112
rect 30009 40103 30067 40109
rect 30009 40069 30021 40103
rect 30055 40100 30067 40103
rect 31294 40100 31300 40112
rect 30055 40072 31300 40100
rect 30055 40069 30067 40072
rect 30009 40063 30067 40069
rect 31294 40060 31300 40072
rect 31352 40060 31358 40112
rect 31726 40100 31754 40128
rect 32217 40103 32275 40109
rect 32217 40100 32229 40103
rect 31726 40072 32229 40100
rect 32217 40069 32229 40072
rect 32263 40069 32275 40103
rect 32217 40063 32275 40069
rect 33137 40103 33195 40109
rect 33137 40069 33149 40103
rect 33183 40069 33195 40103
rect 33137 40063 33195 40069
rect 33237 40103 33295 40109
rect 33237 40069 33249 40103
rect 33283 40100 33295 40103
rect 34514 40100 34520 40112
rect 33283 40072 34520 40100
rect 33283 40069 33295 40072
rect 33237 40063 33295 40069
rect 27893 40035 27951 40041
rect 27893 40032 27905 40035
rect 27672 40004 27905 40032
rect 27672 39992 27678 40004
rect 27893 40001 27905 40004
rect 27939 40001 27951 40035
rect 27893 39995 27951 40001
rect 28169 40035 28227 40041
rect 28169 40001 28181 40035
rect 28215 40001 28227 40035
rect 28169 39995 28227 40001
rect 30374 39992 30380 40044
rect 30432 40032 30438 40044
rect 30653 40035 30711 40041
rect 30653 40032 30665 40035
rect 30432 40004 30665 40032
rect 30432 39992 30438 40004
rect 30653 40001 30665 40004
rect 30699 40001 30711 40035
rect 30834 40032 30840 40044
rect 30795 40004 30840 40032
rect 30653 39995 30711 40001
rect 30834 39992 30840 40004
rect 30892 39992 30898 40044
rect 31021 40035 31079 40041
rect 31021 40001 31033 40035
rect 31067 40032 31079 40035
rect 32122 40032 32128 40044
rect 31067 40004 32128 40032
rect 31067 40001 31079 40004
rect 31021 39995 31079 40001
rect 32122 39992 32128 40004
rect 32180 39992 32186 40044
rect 32306 39992 32312 40044
rect 32364 40032 32370 40044
rect 32766 40032 32772 40044
rect 32364 40004 32772 40032
rect 32364 39992 32370 40004
rect 32766 39992 32772 40004
rect 32824 40032 32830 40044
rect 33042 40041 33048 40044
rect 32861 40035 32919 40041
rect 32861 40032 32873 40035
rect 32824 40004 32873 40032
rect 32824 39992 32830 40004
rect 32861 40001 32873 40004
rect 32907 40001 32919 40035
rect 32861 39995 32919 40001
rect 33009 40035 33048 40041
rect 33009 40001 33021 40035
rect 33009 39995 33048 40001
rect 33042 39992 33048 39995
rect 33100 39992 33106 40044
rect 33152 39976 33180 40063
rect 34514 40060 34520 40072
rect 34572 40060 34578 40112
rect 39482 40100 39488 40112
rect 39443 40072 39488 40100
rect 39482 40060 39488 40072
rect 39540 40060 39546 40112
rect 40310 40100 40316 40112
rect 39776 40072 40316 40100
rect 33326 40035 33384 40041
rect 33326 40032 33338 40035
rect 33244 40004 33338 40032
rect 33244 39976 33272 40004
rect 33326 40001 33338 40004
rect 33372 40001 33384 40035
rect 33326 39995 33384 40001
rect 34701 40035 34759 40041
rect 34701 40001 34713 40035
rect 34747 40032 34759 40035
rect 35434 40032 35440 40044
rect 34747 40004 35440 40032
rect 34747 40001 34759 40004
rect 34701 39995 34759 40001
rect 35434 39992 35440 40004
rect 35492 39992 35498 40044
rect 37737 40035 37795 40041
rect 37737 40001 37749 40035
rect 37783 40032 37795 40035
rect 38378 40032 38384 40044
rect 37783 40004 38384 40032
rect 37783 40001 37795 40004
rect 37737 39995 37795 40001
rect 38378 39992 38384 40004
rect 38436 39992 38442 40044
rect 39776 40041 39804 40072
rect 40310 40060 40316 40072
rect 40368 40060 40374 40112
rect 40586 40100 40592 40112
rect 40547 40072 40592 40100
rect 40586 40060 40592 40072
rect 40644 40060 40650 40112
rect 40773 40103 40831 40109
rect 40773 40069 40785 40103
rect 40819 40100 40831 40103
rect 40819 40072 41736 40100
rect 40819 40069 40831 40072
rect 40773 40063 40831 40069
rect 38565 40035 38623 40041
rect 38565 40001 38577 40035
rect 38611 40001 38623 40035
rect 39669 40035 39727 40041
rect 39669 40032 39681 40035
rect 38565 39995 38623 40001
rect 39500 40004 39681 40032
rect 23658 39964 23664 39976
rect 23619 39936 23664 39964
rect 23658 39924 23664 39936
rect 23716 39924 23722 39976
rect 24397 39967 24455 39973
rect 24397 39933 24409 39967
rect 24443 39933 24455 39967
rect 24397 39927 24455 39933
rect 2222 39788 2228 39840
rect 2280 39828 2286 39840
rect 2409 39831 2467 39837
rect 2409 39828 2421 39831
rect 2280 39800 2421 39828
rect 2280 39788 2286 39800
rect 2409 39797 2421 39800
rect 2455 39797 2467 39831
rect 24412 39828 24440 39927
rect 25406 39924 25412 39976
rect 25464 39964 25470 39976
rect 26329 39967 26387 39973
rect 26329 39964 26341 39967
rect 25464 39936 26341 39964
rect 25464 39924 25470 39936
rect 26329 39933 26341 39936
rect 26375 39933 26387 39967
rect 26329 39927 26387 39933
rect 33134 39924 33140 39976
rect 33192 39924 33198 39976
rect 33226 39924 33232 39976
rect 33284 39924 33290 39976
rect 34882 39964 34888 39976
rect 34843 39936 34888 39964
rect 34882 39924 34888 39936
rect 34940 39924 34946 39976
rect 34974 39924 34980 39976
rect 35032 39964 35038 39976
rect 35032 39936 35077 39964
rect 35032 39924 35038 39936
rect 36814 39924 36820 39976
rect 36872 39964 36878 39976
rect 37553 39967 37611 39973
rect 37553 39964 37565 39967
rect 36872 39936 37565 39964
rect 36872 39924 36878 39936
rect 37553 39933 37565 39936
rect 37599 39964 37611 39967
rect 38580 39964 38608 39995
rect 39500 39976 39528 40004
rect 39669 40001 39681 40004
rect 39715 40001 39727 40035
rect 39669 39995 39727 40001
rect 39761 40035 39819 40041
rect 39761 40001 39773 40035
rect 39807 40001 39819 40035
rect 41506 40032 41512 40044
rect 41467 40004 41512 40032
rect 39761 39995 39819 40001
rect 41506 39992 41512 40004
rect 41564 39992 41570 40044
rect 41708 40041 41736 40072
rect 45554 40060 45560 40112
rect 45612 40100 45618 40112
rect 45830 40100 45836 40112
rect 45612 40072 45836 40100
rect 45612 40060 45618 40072
rect 45830 40060 45836 40072
rect 45888 40100 45894 40112
rect 46658 40100 46664 40112
rect 45888 40072 46664 40100
rect 45888 40060 45894 40072
rect 46658 40060 46664 40072
rect 46716 40060 46722 40112
rect 46845 40103 46903 40109
rect 46845 40069 46857 40103
rect 46891 40100 46903 40103
rect 47118 40100 47124 40112
rect 46891 40072 47124 40100
rect 46891 40069 46903 40072
rect 46845 40063 46903 40069
rect 47118 40060 47124 40072
rect 47176 40060 47182 40112
rect 41693 40035 41751 40041
rect 41693 40001 41705 40035
rect 41739 40032 41751 40035
rect 42242 40032 42248 40044
rect 41739 40004 42248 40032
rect 41739 40001 41751 40004
rect 41693 39995 41751 40001
rect 42242 39992 42248 40004
rect 42300 40032 42306 40044
rect 42702 40032 42708 40044
rect 42300 40004 42708 40032
rect 42300 39992 42306 40004
rect 42702 39992 42708 40004
rect 42760 39992 42766 40044
rect 44085 40035 44143 40041
rect 44085 40001 44097 40035
rect 44131 40032 44143 40035
rect 44818 40032 44824 40044
rect 44131 40004 44824 40032
rect 44131 40001 44143 40004
rect 44085 39995 44143 40001
rect 44818 39992 44824 40004
rect 44876 39992 44882 40044
rect 45097 40035 45155 40041
rect 45097 40001 45109 40035
rect 45143 40032 45155 40035
rect 46566 40032 46572 40044
rect 45143 40004 46572 40032
rect 45143 40001 45155 40004
rect 45097 39995 45155 40001
rect 37599 39936 38608 39964
rect 37599 39933 37611 39936
rect 37553 39927 37611 39933
rect 39482 39924 39488 39976
rect 39540 39924 39546 39976
rect 39850 39924 39856 39976
rect 39908 39964 39914 39976
rect 45112 39964 45140 39995
rect 46566 39992 46572 40004
rect 46624 40032 46630 40044
rect 48056 40041 48084 40140
rect 48866 40128 48872 40140
rect 48924 40128 48930 40180
rect 49160 40140 50108 40168
rect 48774 40060 48780 40112
rect 48832 40100 48838 40112
rect 49160 40100 49188 40140
rect 48832 40072 49188 40100
rect 48832 40060 48838 40072
rect 49234 40060 49240 40112
rect 49292 40100 49298 40112
rect 49292 40072 49337 40100
rect 49292 40060 49298 40072
rect 48041 40035 48099 40041
rect 46624 40004 46934 40032
rect 46624 39992 46630 40004
rect 39908 39936 45140 39964
rect 45189 39967 45247 39973
rect 39908 39924 39914 39936
rect 45189 39933 45201 39967
rect 45235 39964 45247 39967
rect 45554 39964 45560 39976
rect 45235 39936 45560 39964
rect 45235 39933 45247 39936
rect 45189 39927 45247 39933
rect 45554 39924 45560 39936
rect 45612 39924 45618 39976
rect 46906 39964 46934 40004
rect 48041 40001 48053 40035
rect 48087 40001 48099 40035
rect 48041 39995 48099 40001
rect 49878 39992 49884 40044
rect 49936 40032 49942 40044
rect 50080 40041 50108 40140
rect 51074 40128 51080 40180
rect 51132 40168 51138 40180
rect 51445 40171 51503 40177
rect 51445 40168 51457 40171
rect 51132 40140 51457 40168
rect 51132 40128 51138 40140
rect 51445 40137 51457 40140
rect 51491 40137 51503 40171
rect 51445 40131 51503 40137
rect 51629 40171 51687 40177
rect 51629 40137 51641 40171
rect 51675 40168 51687 40171
rect 52730 40168 52736 40180
rect 51675 40140 52736 40168
rect 51675 40137 51687 40140
rect 51629 40131 51687 40137
rect 52730 40128 52736 40140
rect 52788 40128 52794 40180
rect 52822 40128 52828 40180
rect 52880 40168 52886 40180
rect 56226 40168 56232 40180
rect 52880 40140 56232 40168
rect 52880 40128 52886 40140
rect 51261 40103 51319 40109
rect 51261 40069 51273 40103
rect 51307 40100 51319 40103
rect 51307 40072 51764 40100
rect 51307 40069 51319 40072
rect 51261 40063 51319 40069
rect 51736 40044 51764 40072
rect 50065 40035 50123 40041
rect 49936 40004 49981 40032
rect 49936 39992 49942 40004
rect 50065 40001 50077 40035
rect 50111 40001 50123 40035
rect 50065 39995 50123 40001
rect 50617 40035 50675 40041
rect 50617 40001 50629 40035
rect 50663 40001 50675 40035
rect 50798 40032 50804 40044
rect 50759 40004 50804 40032
rect 50617 39995 50675 40001
rect 48225 39967 48283 39973
rect 48225 39964 48237 39967
rect 46906 39936 48237 39964
rect 48225 39933 48237 39936
rect 48271 39933 48283 39967
rect 50632 39964 50660 39995
rect 50798 39992 50804 40004
rect 50856 39992 50862 40044
rect 51166 39992 51172 40044
rect 51224 40032 51230 40044
rect 51537 40035 51595 40041
rect 51537 40032 51549 40035
rect 51224 40004 51549 40032
rect 51224 39992 51230 40004
rect 51537 40001 51549 40004
rect 51583 40001 51595 40035
rect 51537 39995 51595 40001
rect 51718 39992 51724 40044
rect 51776 39992 51782 40044
rect 51902 39992 51908 40044
rect 51960 40032 51966 40044
rect 53944 40041 53972 40140
rect 56226 40128 56232 40140
rect 56284 40128 56290 40180
rect 56410 40128 56416 40180
rect 56468 40168 56474 40180
rect 56505 40171 56563 40177
rect 56505 40168 56517 40171
rect 56468 40140 56517 40168
rect 56468 40128 56474 40140
rect 56505 40137 56517 40140
rect 56551 40137 56563 40171
rect 56505 40131 56563 40137
rect 54021 40103 54079 40109
rect 54021 40069 54033 40103
rect 54067 40100 54079 40103
rect 55766 40100 55772 40112
rect 54067 40072 54800 40100
rect 54067 40069 54079 40072
rect 54021 40063 54079 40069
rect 54772 40044 54800 40072
rect 55232 40072 55772 40100
rect 55232 40044 55260 40072
rect 55766 40060 55772 40072
rect 55824 40060 55830 40112
rect 52917 40035 52975 40041
rect 51960 40030 52868 40032
rect 52917 40030 52929 40035
rect 51960 40004 52929 40030
rect 51960 39992 51966 40004
rect 52840 40002 52929 40004
rect 52917 40001 52929 40002
rect 52963 40001 52975 40035
rect 52917 39995 52975 40001
rect 53929 40035 53987 40041
rect 53929 40001 53941 40035
rect 53975 40001 53987 40035
rect 54110 40032 54116 40044
rect 54071 40004 54116 40032
rect 53929 39995 53987 40001
rect 54110 39992 54116 40004
rect 54168 39992 54174 40044
rect 54754 40032 54760 40044
rect 54715 40004 54760 40032
rect 54754 39992 54760 40004
rect 54812 39992 54818 40044
rect 55214 40032 55220 40044
rect 54864 40004 55220 40032
rect 51350 39964 51356 39976
rect 50632 39936 51356 39964
rect 48225 39927 48283 39933
rect 51350 39924 51356 39936
rect 51408 39924 51414 39976
rect 54864 39973 54892 40004
rect 55214 39992 55220 40004
rect 55272 39992 55278 40044
rect 55306 39992 55312 40044
rect 55364 40032 55370 40044
rect 56137 40035 56195 40041
rect 56137 40032 56149 40035
rect 55364 40004 56149 40032
rect 55364 39992 55370 40004
rect 56137 40001 56149 40004
rect 56183 40032 56195 40035
rect 56318 40032 56324 40044
rect 56183 40004 56324 40032
rect 56183 40001 56195 40004
rect 56137 39995 56195 40001
rect 56318 39992 56324 40004
rect 56376 39992 56382 40044
rect 57882 40032 57888 40044
rect 57843 40004 57888 40032
rect 57882 39992 57888 40004
rect 57940 39992 57946 40044
rect 53009 39967 53067 39973
rect 53009 39964 53021 39967
rect 51736 39936 53021 39964
rect 28902 39896 28908 39908
rect 28863 39868 28908 39896
rect 28902 39856 28908 39868
rect 28960 39856 28966 39908
rect 30282 39856 30288 39908
rect 30340 39896 30346 39908
rect 48314 39896 48320 39908
rect 30340 39868 48320 39896
rect 30340 39856 30346 39868
rect 48314 39856 48320 39868
rect 48372 39856 48378 39908
rect 50709 39899 50767 39905
rect 49160 39868 49464 39896
rect 27522 39828 27528 39840
rect 24412 39800 27528 39828
rect 2409 39791 2467 39797
rect 27522 39788 27528 39800
rect 27580 39828 27586 39840
rect 28994 39828 29000 39840
rect 27580 39800 29000 39828
rect 27580 39788 27586 39800
rect 28994 39788 29000 39800
rect 29052 39788 29058 39840
rect 31846 39788 31852 39840
rect 31904 39828 31910 39840
rect 32309 39831 32367 39837
rect 32309 39828 32321 39831
rect 31904 39800 32321 39828
rect 31904 39788 31910 39800
rect 32309 39797 32321 39800
rect 32355 39828 32367 39831
rect 32582 39828 32588 39840
rect 32355 39800 32588 39828
rect 32355 39797 32367 39800
rect 32309 39791 32367 39797
rect 32582 39788 32588 39800
rect 32640 39788 32646 39840
rect 33226 39788 33232 39840
rect 33284 39828 33290 39840
rect 33505 39831 33563 39837
rect 33505 39828 33517 39831
rect 33284 39800 33517 39828
rect 33284 39788 33290 39800
rect 33505 39797 33517 39800
rect 33551 39797 33563 39831
rect 34514 39828 34520 39840
rect 34475 39800 34520 39828
rect 33505 39791 33563 39797
rect 34514 39788 34520 39800
rect 34572 39788 34578 39840
rect 39485 39831 39543 39837
rect 39485 39797 39497 39831
rect 39531 39828 39543 39831
rect 40126 39828 40132 39840
rect 39531 39800 40132 39828
rect 39531 39797 39543 39800
rect 39485 39791 39543 39797
rect 40126 39788 40132 39800
rect 40184 39788 40190 39840
rect 41414 39788 41420 39840
rect 41472 39828 41478 39840
rect 41509 39831 41567 39837
rect 41509 39828 41521 39831
rect 41472 39800 41521 39828
rect 41472 39788 41478 39800
rect 41509 39797 41521 39800
rect 41555 39797 41567 39831
rect 41509 39791 41567 39797
rect 44174 39788 44180 39840
rect 44232 39828 44238 39840
rect 44269 39831 44327 39837
rect 44269 39828 44281 39831
rect 44232 39800 44281 39828
rect 44232 39788 44238 39800
rect 44269 39797 44281 39800
rect 44315 39797 44327 39831
rect 44269 39791 44327 39797
rect 44358 39788 44364 39840
rect 44416 39828 44422 39840
rect 45094 39828 45100 39840
rect 44416 39800 45100 39828
rect 44416 39788 44422 39800
rect 45094 39788 45100 39800
rect 45152 39788 45158 39840
rect 45370 39828 45376 39840
rect 45331 39800 45376 39828
rect 45370 39788 45376 39800
rect 45428 39788 45434 39840
rect 45554 39788 45560 39840
rect 45612 39828 45618 39840
rect 46474 39828 46480 39840
rect 45612 39800 46480 39828
rect 45612 39788 45618 39800
rect 46474 39788 46480 39800
rect 46532 39828 46538 39840
rect 46937 39831 46995 39837
rect 46937 39828 46949 39831
rect 46532 39800 46949 39828
rect 46532 39788 46538 39800
rect 46937 39797 46949 39800
rect 46983 39797 46995 39831
rect 46937 39791 46995 39797
rect 47486 39788 47492 39840
rect 47544 39828 47550 39840
rect 49160 39828 49188 39868
rect 49326 39828 49332 39840
rect 47544 39800 49188 39828
rect 49287 39800 49332 39828
rect 47544 39788 47550 39800
rect 49326 39788 49332 39800
rect 49384 39788 49390 39840
rect 49436 39828 49464 39868
rect 50709 39865 50721 39899
rect 50755 39896 50767 39899
rect 51736 39896 51764 39936
rect 53009 39933 53021 39936
rect 53055 39933 53067 39967
rect 53009 39927 53067 39933
rect 54849 39967 54907 39973
rect 54849 39933 54861 39967
rect 54895 39933 54907 39967
rect 55122 39964 55128 39976
rect 55083 39936 55128 39964
rect 54849 39927 54907 39933
rect 55122 39924 55128 39936
rect 55180 39924 55186 39976
rect 56229 39967 56287 39973
rect 56229 39933 56241 39967
rect 56275 39964 56287 39967
rect 56410 39964 56416 39976
rect 56275 39936 56416 39964
rect 56275 39933 56287 39936
rect 56229 39927 56287 39933
rect 56410 39924 56416 39936
rect 56468 39924 56474 39976
rect 50755 39868 51764 39896
rect 51813 39899 51871 39905
rect 50755 39865 50767 39868
rect 50709 39859 50767 39865
rect 51813 39865 51825 39899
rect 51859 39896 51871 39899
rect 52822 39896 52828 39908
rect 51859 39868 52828 39896
rect 51859 39865 51871 39868
rect 51813 39859 51871 39865
rect 52822 39856 52828 39868
rect 52880 39856 52886 39908
rect 53926 39856 53932 39908
rect 53984 39896 53990 39908
rect 58069 39899 58127 39905
rect 58069 39896 58081 39899
rect 53984 39868 58081 39896
rect 53984 39856 53990 39868
rect 58069 39865 58081 39868
rect 58115 39865 58127 39899
rect 58069 39859 58127 39865
rect 49973 39831 50031 39837
rect 49973 39828 49985 39831
rect 49436 39800 49985 39828
rect 49973 39797 49985 39800
rect 50019 39797 50031 39831
rect 53190 39828 53196 39840
rect 53151 39800 53196 39828
rect 49973 39791 50031 39797
rect 53190 39788 53196 39800
rect 53248 39788 53254 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 22833 39627 22891 39633
rect 22833 39593 22845 39627
rect 22879 39624 22891 39627
rect 24302 39624 24308 39636
rect 22879 39596 24308 39624
rect 22879 39593 22891 39596
rect 22833 39587 22891 39593
rect 24302 39584 24308 39596
rect 24360 39584 24366 39636
rect 24397 39627 24455 39633
rect 24397 39593 24409 39627
rect 24443 39624 24455 39627
rect 24486 39624 24492 39636
rect 24443 39596 24492 39624
rect 24443 39593 24455 39596
rect 24397 39587 24455 39593
rect 24486 39584 24492 39596
rect 24544 39584 24550 39636
rect 24578 39584 24584 39636
rect 24636 39624 24642 39636
rect 25685 39627 25743 39633
rect 25685 39624 25697 39627
rect 24636 39596 25697 39624
rect 24636 39584 24642 39596
rect 25685 39593 25697 39596
rect 25731 39624 25743 39627
rect 33042 39624 33048 39636
rect 25731 39596 33048 39624
rect 25731 39593 25743 39596
rect 25685 39587 25743 39593
rect 33042 39584 33048 39596
rect 33100 39624 33106 39636
rect 33100 39596 35296 39624
rect 33100 39584 33106 39596
rect 23934 39516 23940 39568
rect 23992 39556 23998 39568
rect 28997 39559 29055 39565
rect 23992 39528 24256 39556
rect 23992 39516 23998 39528
rect 21910 39488 21916 39500
rect 21100 39460 21916 39488
rect 3789 39423 3847 39429
rect 3789 39389 3801 39423
rect 3835 39420 3847 39423
rect 3878 39420 3884 39432
rect 3835 39392 3884 39420
rect 3835 39389 3847 39392
rect 3789 39383 3847 39389
rect 3878 39380 3884 39392
rect 3936 39420 3942 39432
rect 4614 39420 4620 39432
rect 3936 39392 4620 39420
rect 3936 39380 3942 39392
rect 4614 39380 4620 39392
rect 4672 39380 4678 39432
rect 20898 39420 20904 39432
rect 20859 39392 20904 39420
rect 20898 39380 20904 39392
rect 20956 39380 20962 39432
rect 21100 39429 21128 39460
rect 21910 39448 21916 39460
rect 21968 39488 21974 39500
rect 23845 39491 23903 39497
rect 23845 39488 23857 39491
rect 21968 39460 23857 39488
rect 21968 39448 21974 39460
rect 23845 39457 23857 39460
rect 23891 39488 23903 39491
rect 24118 39488 24124 39500
rect 23891 39460 24124 39488
rect 23891 39457 23903 39460
rect 23845 39451 23903 39457
rect 24118 39448 24124 39460
rect 24176 39448 24182 39500
rect 24228 39488 24256 39528
rect 24596 39528 24808 39556
rect 24596 39488 24624 39528
rect 24228 39460 24624 39488
rect 21085 39423 21143 39429
rect 21085 39389 21097 39423
rect 21131 39389 21143 39423
rect 22738 39420 22744 39432
rect 22699 39392 22744 39420
rect 21085 39383 21143 39389
rect 22738 39380 22744 39392
rect 22796 39380 22802 39432
rect 22925 39423 22983 39429
rect 22925 39389 22937 39423
rect 22971 39420 22983 39423
rect 24578 39420 24584 39432
rect 22971 39392 24584 39420
rect 22971 39389 22983 39392
rect 22925 39383 22983 39389
rect 24578 39380 24584 39392
rect 24636 39429 24642 39432
rect 24780 39429 24808 39528
rect 28997 39525 29009 39559
rect 29043 39556 29055 39559
rect 29822 39556 29828 39568
rect 29043 39528 29828 39556
rect 29043 39525 29055 39528
rect 28997 39519 29055 39525
rect 29822 39516 29828 39528
rect 29880 39516 29886 39568
rect 32122 39516 32128 39568
rect 32180 39556 32186 39568
rect 33686 39556 33692 39568
rect 32180 39528 33692 39556
rect 32180 39516 32186 39528
rect 33686 39516 33692 39528
rect 33744 39516 33750 39568
rect 28902 39448 28908 39500
rect 28960 39488 28966 39500
rect 28960 39460 34459 39488
rect 28960 39448 28966 39460
rect 24636 39423 24685 39429
rect 24636 39389 24639 39423
rect 24673 39389 24685 39423
rect 24636 39383 24685 39389
rect 24765 39423 24823 39429
rect 24765 39389 24777 39423
rect 24811 39389 24823 39423
rect 24765 39383 24823 39389
rect 24636 39380 24642 39383
rect 24854 39380 24860 39432
rect 24912 39429 24918 39432
rect 24912 39420 24920 39429
rect 24912 39392 24957 39420
rect 24912 39383 24920 39392
rect 24912 39380 24918 39383
rect 25038 39380 25044 39432
rect 25096 39420 25102 39432
rect 25096 39392 25141 39420
rect 25096 39380 25102 39392
rect 25498 39380 25504 39432
rect 25556 39420 25562 39432
rect 25593 39423 25651 39429
rect 25593 39420 25605 39423
rect 25556 39392 25605 39420
rect 25556 39380 25562 39392
rect 25593 39389 25605 39392
rect 25639 39389 25651 39423
rect 25593 39383 25651 39389
rect 27522 39380 27528 39432
rect 27580 39420 27586 39432
rect 27890 39429 27896 39432
rect 27617 39423 27675 39429
rect 27617 39420 27629 39423
rect 27580 39392 27629 39420
rect 27580 39380 27586 39392
rect 27617 39389 27629 39392
rect 27663 39389 27675 39423
rect 27884 39420 27896 39429
rect 27851 39392 27896 39420
rect 27617 39383 27675 39389
rect 27884 39383 27896 39392
rect 27890 39380 27896 39383
rect 27948 39380 27954 39432
rect 29917 39423 29975 39429
rect 29917 39389 29929 39423
rect 29963 39420 29975 39423
rect 30190 39420 30196 39432
rect 29963 39392 30196 39420
rect 29963 39389 29975 39392
rect 29917 39383 29975 39389
rect 30190 39380 30196 39392
rect 30248 39380 30254 39432
rect 30745 39423 30803 39429
rect 30745 39389 30757 39423
rect 30791 39420 30803 39423
rect 31478 39420 31484 39432
rect 30791 39392 31484 39420
rect 30791 39389 30803 39392
rect 30745 39383 30803 39389
rect 31478 39380 31484 39392
rect 31536 39380 31542 39432
rect 31754 39420 31760 39432
rect 31726 39380 31760 39420
rect 31812 39420 31818 39432
rect 31905 39423 31963 39429
rect 31812 39392 31857 39420
rect 31812 39380 31818 39392
rect 31905 39389 31917 39423
rect 31951 39420 31963 39423
rect 32122 39420 32128 39432
rect 31951 39389 31984 39420
rect 32083 39392 32128 39420
rect 31905 39383 31984 39389
rect 23661 39355 23719 39361
rect 23661 39321 23673 39355
rect 23707 39352 23719 39355
rect 23842 39352 23848 39364
rect 23707 39324 23848 39352
rect 23707 39321 23719 39324
rect 23661 39315 23719 39321
rect 23842 39312 23848 39324
rect 23900 39312 23906 39364
rect 30837 39355 30895 39361
rect 30837 39352 30849 39355
rect 28920 39324 30849 39352
rect 2406 39244 2412 39296
rect 2464 39284 2470 39296
rect 3881 39287 3939 39293
rect 3881 39284 3893 39287
rect 2464 39256 3893 39284
rect 2464 39244 2470 39256
rect 3881 39253 3893 39256
rect 3927 39253 3939 39287
rect 21082 39284 21088 39296
rect 21043 39256 21088 39284
rect 3881 39247 3939 39253
rect 21082 39244 21088 39256
rect 21140 39244 21146 39296
rect 27614 39244 27620 39296
rect 27672 39284 27678 39296
rect 28920 39284 28948 39324
rect 30837 39321 30849 39324
rect 30883 39352 30895 39355
rect 31726 39352 31754 39380
rect 30883 39324 31754 39352
rect 30883 39321 30895 39324
rect 30837 39315 30895 39321
rect 27672 39256 28948 39284
rect 30009 39287 30067 39293
rect 27672 39244 27678 39256
rect 30009 39253 30021 39287
rect 30055 39284 30067 39287
rect 30282 39284 30288 39296
rect 30055 39256 30288 39284
rect 30055 39253 30067 39256
rect 30009 39247 30067 39253
rect 30282 39244 30288 39256
rect 30340 39244 30346 39296
rect 31956 39284 31984 39383
rect 32122 39380 32128 39392
rect 32180 39380 32186 39432
rect 32263 39423 32321 39429
rect 32263 39389 32275 39423
rect 32309 39420 32321 39423
rect 32490 39420 32496 39432
rect 32309 39392 32496 39420
rect 32309 39389 32321 39392
rect 32263 39383 32321 39389
rect 32490 39380 32496 39392
rect 32548 39420 32554 39432
rect 32548 39392 32720 39420
rect 32548 39380 32554 39392
rect 32033 39355 32091 39361
rect 32033 39321 32045 39355
rect 32079 39352 32091 39355
rect 32582 39352 32588 39364
rect 32079 39324 32588 39352
rect 32079 39321 32091 39324
rect 32033 39315 32091 39321
rect 32582 39312 32588 39324
rect 32640 39312 32646 39364
rect 32214 39284 32220 39296
rect 31956 39256 32220 39284
rect 32214 39244 32220 39256
rect 32272 39244 32278 39296
rect 32398 39284 32404 39296
rect 32359 39256 32404 39284
rect 32398 39244 32404 39256
rect 32456 39244 32462 39296
rect 32692 39284 32720 39392
rect 32766 39380 32772 39432
rect 32824 39420 32830 39432
rect 33024 39429 33052 39460
rect 32861 39423 32919 39429
rect 32861 39420 32873 39423
rect 32824 39392 32873 39420
rect 32824 39380 32830 39392
rect 32861 39389 32873 39392
rect 32907 39389 32919 39423
rect 32861 39383 32919 39389
rect 33009 39423 33067 39429
rect 33009 39389 33021 39423
rect 33055 39389 33067 39423
rect 33134 39420 33140 39432
rect 33095 39392 33140 39420
rect 33009 39383 33067 39389
rect 33134 39380 33140 39392
rect 33192 39380 33198 39432
rect 33318 39380 33324 39432
rect 33376 39429 33382 39432
rect 33376 39423 33403 39429
rect 33391 39389 33403 39423
rect 33376 39383 33403 39389
rect 33376 39380 33382 39383
rect 33229 39355 33287 39361
rect 33229 39321 33241 39355
rect 33275 39352 33287 39355
rect 34330 39352 34336 39364
rect 33275 39324 34336 39352
rect 33275 39321 33287 39324
rect 33229 39315 33287 39321
rect 34330 39312 34336 39324
rect 34388 39312 34394 39364
rect 34431 39352 34459 39460
rect 34790 39448 34796 39500
rect 34848 39488 34854 39500
rect 35161 39491 35219 39497
rect 35161 39488 35173 39491
rect 34848 39460 35173 39488
rect 34848 39448 34854 39460
rect 35161 39457 35173 39460
rect 35207 39457 35219 39491
rect 35161 39451 35219 39457
rect 34882 39420 34888 39432
rect 34843 39392 34888 39420
rect 34882 39380 34888 39392
rect 34940 39380 34946 39432
rect 34977 39423 35035 39429
rect 34977 39389 34989 39423
rect 35023 39389 35035 39423
rect 34977 39383 35035 39389
rect 35069 39423 35127 39429
rect 35069 39389 35081 39423
rect 35115 39420 35127 39423
rect 35268 39420 35296 39596
rect 39574 39584 39580 39636
rect 39632 39624 39638 39636
rect 39853 39627 39911 39633
rect 39853 39624 39865 39627
rect 39632 39596 39865 39624
rect 39632 39584 39638 39596
rect 39853 39593 39865 39596
rect 39899 39624 39911 39627
rect 40126 39624 40132 39636
rect 39899 39596 40132 39624
rect 39899 39593 39911 39596
rect 39853 39587 39911 39593
rect 40126 39584 40132 39596
rect 40184 39584 40190 39636
rect 40313 39627 40371 39633
rect 40313 39593 40325 39627
rect 40359 39624 40371 39627
rect 40954 39624 40960 39636
rect 40359 39596 40960 39624
rect 40359 39593 40371 39596
rect 40313 39587 40371 39593
rect 40954 39584 40960 39596
rect 41012 39584 41018 39636
rect 41598 39584 41604 39636
rect 41656 39624 41662 39636
rect 41874 39624 41880 39636
rect 41656 39596 41880 39624
rect 41656 39584 41662 39596
rect 41874 39584 41880 39596
rect 41932 39624 41938 39636
rect 44358 39624 44364 39636
rect 41932 39596 44364 39624
rect 41932 39584 41938 39596
rect 44358 39584 44364 39596
rect 44416 39584 44422 39636
rect 45186 39624 45192 39636
rect 44928 39596 45192 39624
rect 35434 39516 35440 39568
rect 35492 39556 35498 39568
rect 44928 39556 44956 39596
rect 45186 39584 45192 39596
rect 45244 39584 45250 39636
rect 45278 39584 45284 39636
rect 45336 39624 45342 39636
rect 47210 39624 47216 39636
rect 45336 39596 47216 39624
rect 45336 39584 45342 39596
rect 47210 39584 47216 39596
rect 47268 39584 47274 39636
rect 48409 39627 48467 39633
rect 48409 39593 48421 39627
rect 48455 39624 48467 39627
rect 54110 39624 54116 39636
rect 48455 39596 54116 39624
rect 48455 39593 48467 39596
rect 48409 39587 48467 39593
rect 54110 39584 54116 39596
rect 54168 39584 54174 39636
rect 55490 39584 55496 39636
rect 55548 39624 55554 39636
rect 55769 39627 55827 39633
rect 55769 39624 55781 39627
rect 55548 39596 55781 39624
rect 55548 39584 55554 39596
rect 55769 39593 55781 39596
rect 55815 39593 55827 39627
rect 56410 39624 56416 39636
rect 56371 39596 56416 39624
rect 55769 39587 55827 39593
rect 56410 39584 56416 39596
rect 56468 39584 56474 39636
rect 56778 39624 56784 39636
rect 56739 39596 56784 39624
rect 56778 39584 56784 39596
rect 56836 39584 56842 39636
rect 35492 39528 44956 39556
rect 35492 39516 35498 39528
rect 45002 39516 45008 39568
rect 45060 39556 45066 39568
rect 45554 39556 45560 39568
rect 45060 39528 45560 39556
rect 45060 39516 45066 39528
rect 45554 39516 45560 39528
rect 45612 39516 45618 39568
rect 46658 39516 46664 39568
rect 46716 39556 46722 39568
rect 49326 39556 49332 39568
rect 46716 39528 49332 39556
rect 46716 39516 46722 39528
rect 49326 39516 49332 39528
rect 49384 39516 49390 39568
rect 54757 39559 54815 39565
rect 54757 39525 54769 39559
rect 54803 39556 54815 39559
rect 55214 39556 55220 39568
rect 54803 39528 55220 39556
rect 54803 39525 54815 39528
rect 54757 39519 54815 39525
rect 55214 39516 55220 39528
rect 55272 39516 55278 39568
rect 55585 39559 55643 39565
rect 55585 39525 55597 39559
rect 55631 39525 55643 39559
rect 55585 39519 55643 39525
rect 38654 39448 38660 39500
rect 38712 39488 38718 39500
rect 39945 39491 40003 39497
rect 39945 39488 39957 39491
rect 38712 39460 39957 39488
rect 38712 39448 38718 39460
rect 39945 39457 39957 39460
rect 39991 39457 40003 39491
rect 39945 39451 40003 39457
rect 40402 39448 40408 39500
rect 40460 39488 40466 39500
rect 41049 39491 41107 39497
rect 41049 39488 41061 39491
rect 40460 39460 41061 39488
rect 40460 39448 40466 39460
rect 41049 39457 41061 39460
rect 41095 39457 41107 39491
rect 41049 39451 41107 39457
rect 44453 39491 44511 39497
rect 44453 39457 44465 39491
rect 44499 39488 44511 39491
rect 48869 39491 48927 39497
rect 48869 39488 48881 39491
rect 44499 39460 45508 39488
rect 44499 39457 44511 39460
rect 44453 39451 44511 39457
rect 37274 39420 37280 39432
rect 35115 39392 37280 39420
rect 35115 39389 35127 39392
rect 35069 39383 35127 39389
rect 34992 39352 35020 39383
rect 37274 39380 37280 39392
rect 37332 39380 37338 39432
rect 39298 39380 39304 39432
rect 39356 39420 39362 39432
rect 40034 39420 40040 39432
rect 39356 39392 40040 39420
rect 39356 39380 39362 39392
rect 40034 39380 40040 39392
rect 40092 39420 40098 39432
rect 40129 39423 40187 39429
rect 40129 39420 40141 39423
rect 40092 39392 40141 39420
rect 40092 39380 40098 39392
rect 40129 39389 40141 39392
rect 40175 39389 40187 39423
rect 40129 39383 40187 39389
rect 40218 39380 40224 39432
rect 40276 39420 40282 39432
rect 44269 39423 44327 39429
rect 44269 39420 44281 39423
rect 40276 39392 44281 39420
rect 40276 39380 40282 39392
rect 44269 39389 44281 39392
rect 44315 39420 44327 39423
rect 45002 39420 45008 39432
rect 44315 39392 45008 39420
rect 44315 39389 44327 39392
rect 44269 39383 44327 39389
rect 45002 39380 45008 39392
rect 45060 39380 45066 39432
rect 45278 39420 45284 39432
rect 45239 39392 45284 39420
rect 45278 39380 45284 39392
rect 45336 39380 45342 39432
rect 45480 39429 45508 39460
rect 45756 39460 48881 39488
rect 45373 39423 45431 39429
rect 45373 39389 45385 39423
rect 45419 39389 45431 39423
rect 45373 39383 45431 39389
rect 45465 39423 45523 39429
rect 45465 39389 45477 39423
rect 45511 39389 45523 39423
rect 45646 39420 45652 39432
rect 45607 39392 45652 39420
rect 45465 39383 45523 39389
rect 35802 39352 35808 39364
rect 34431 39324 34836 39352
rect 34992 39324 35808 39352
rect 33318 39284 33324 39296
rect 32692 39256 33324 39284
rect 33318 39244 33324 39256
rect 33376 39244 33382 39296
rect 33502 39284 33508 39296
rect 33463 39256 33508 39284
rect 33502 39244 33508 39256
rect 33560 39244 33566 39296
rect 34606 39244 34612 39296
rect 34664 39284 34670 39296
rect 34701 39287 34759 39293
rect 34701 39284 34713 39287
rect 34664 39256 34713 39284
rect 34664 39244 34670 39256
rect 34701 39253 34713 39256
rect 34747 39253 34759 39287
rect 34808 39284 34836 39324
rect 35802 39312 35808 39324
rect 35860 39312 35866 39364
rect 39853 39355 39911 39361
rect 39853 39321 39865 39355
rect 39899 39352 39911 39355
rect 39942 39352 39948 39364
rect 39899 39324 39948 39352
rect 39899 39321 39911 39324
rect 39853 39315 39911 39321
rect 39942 39312 39948 39324
rect 40000 39352 40006 39364
rect 40586 39352 40592 39364
rect 40000 39324 40592 39352
rect 40000 39312 40006 39324
rect 40586 39312 40592 39324
rect 40644 39312 40650 39364
rect 40862 39312 40868 39364
rect 40920 39352 40926 39364
rect 44082 39352 44088 39364
rect 40920 39324 40965 39352
rect 44043 39324 44088 39352
rect 40920 39312 40926 39324
rect 44082 39312 44088 39324
rect 44140 39312 44146 39364
rect 44818 39312 44824 39364
rect 44876 39352 44882 39364
rect 45186 39352 45192 39364
rect 44876 39324 45192 39352
rect 44876 39312 44882 39324
rect 45186 39312 45192 39324
rect 45244 39352 45250 39364
rect 45388 39352 45416 39383
rect 45646 39380 45652 39392
rect 45704 39380 45710 39432
rect 45244 39324 45416 39352
rect 45244 39312 45250 39324
rect 35986 39284 35992 39296
rect 34808 39256 35992 39284
rect 34701 39247 34759 39253
rect 35986 39244 35992 39256
rect 36044 39244 36050 39296
rect 37366 39244 37372 39296
rect 37424 39284 37430 39296
rect 37734 39284 37740 39296
rect 37424 39256 37740 39284
rect 37424 39244 37430 39256
rect 37734 39244 37740 39256
rect 37792 39284 37798 39296
rect 38562 39284 38568 39296
rect 37792 39256 38568 39284
rect 37792 39244 37798 39256
rect 38562 39244 38568 39256
rect 38620 39244 38626 39296
rect 44726 39244 44732 39296
rect 44784 39284 44790 39296
rect 45005 39287 45063 39293
rect 45005 39284 45017 39287
rect 44784 39256 45017 39284
rect 44784 39244 44790 39256
rect 45005 39253 45017 39256
rect 45051 39253 45063 39287
rect 45005 39247 45063 39253
rect 45094 39244 45100 39296
rect 45152 39284 45158 39296
rect 45756 39284 45784 39460
rect 48869 39457 48881 39460
rect 48915 39457 48927 39491
rect 51166 39488 51172 39500
rect 51127 39460 51172 39488
rect 48869 39451 48927 39457
rect 51166 39448 51172 39460
rect 51224 39448 51230 39500
rect 54478 39488 54484 39500
rect 54439 39460 54484 39488
rect 54478 39448 54484 39460
rect 54536 39488 54542 39500
rect 55600 39488 55628 39519
rect 54536 39460 55628 39488
rect 54536 39448 54542 39460
rect 48590 39420 48596 39432
rect 48551 39392 48596 39420
rect 48590 39380 48596 39392
rect 48648 39380 48654 39432
rect 48682 39380 48688 39432
rect 48740 39420 48746 39432
rect 48958 39420 48964 39432
rect 48740 39392 48785 39420
rect 48919 39392 48964 39420
rect 48740 39380 48746 39392
rect 48958 39380 48964 39392
rect 49016 39420 49022 39432
rect 50157 39423 50215 39429
rect 50157 39420 50169 39423
rect 49016 39392 50169 39420
rect 49016 39380 49022 39392
rect 50157 39389 50169 39392
rect 50203 39389 50215 39423
rect 50157 39383 50215 39389
rect 50893 39423 50951 39429
rect 50893 39389 50905 39423
rect 50939 39420 50951 39423
rect 51626 39420 51632 39432
rect 50939 39392 51632 39420
rect 50939 39389 50951 39392
rect 50893 39383 50951 39389
rect 51626 39380 51632 39392
rect 51684 39380 51690 39432
rect 53650 39380 53656 39432
rect 53708 39420 53714 39432
rect 54389 39423 54447 39429
rect 54389 39420 54401 39423
rect 53708 39392 54401 39420
rect 53708 39380 53714 39392
rect 54389 39389 54401 39392
rect 54435 39420 54447 39423
rect 55309 39423 55367 39429
rect 55309 39420 55321 39423
rect 54435 39392 55321 39420
rect 54435 39389 54447 39392
rect 54389 39383 54447 39389
rect 55309 39389 55321 39392
rect 55355 39389 55367 39423
rect 56318 39420 56324 39432
rect 56279 39392 56324 39420
rect 55309 39383 55367 39389
rect 56318 39380 56324 39392
rect 56376 39380 56382 39432
rect 57241 39423 57299 39429
rect 57241 39389 57253 39423
rect 57287 39420 57299 39423
rect 57790 39420 57796 39432
rect 57287 39392 57796 39420
rect 57287 39389 57299 39392
rect 57241 39383 57299 39389
rect 57790 39380 57796 39392
rect 57848 39380 57854 39432
rect 48608 39352 48636 39380
rect 50062 39352 50068 39364
rect 48608 39324 50068 39352
rect 50062 39312 50068 39324
rect 50120 39312 50126 39364
rect 45152 39256 45784 39284
rect 45152 39244 45158 39256
rect 47210 39244 47216 39296
rect 47268 39284 47274 39296
rect 49418 39284 49424 39296
rect 47268 39256 49424 39284
rect 47268 39244 47274 39256
rect 49418 39244 49424 39256
rect 49476 39284 49482 39296
rect 50341 39287 50399 39293
rect 50341 39284 50353 39287
rect 49476 39256 50353 39284
rect 49476 39244 49482 39256
rect 50341 39253 50353 39256
rect 50387 39253 50399 39287
rect 50341 39247 50399 39253
rect 50798 39244 50804 39296
rect 50856 39284 50862 39296
rect 51166 39284 51172 39296
rect 50856 39256 51172 39284
rect 50856 39244 50862 39256
rect 51166 39244 51172 39256
rect 51224 39244 51230 39296
rect 57330 39284 57336 39296
rect 57291 39256 57336 39284
rect 57330 39244 57336 39256
rect 57388 39244 57394 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 23382 39040 23388 39092
rect 23440 39080 23446 39092
rect 28902 39080 28908 39092
rect 23440 39052 28908 39080
rect 23440 39040 23446 39052
rect 28902 39040 28908 39052
rect 28960 39040 28966 39092
rect 28997 39083 29055 39089
rect 28997 39049 29009 39083
rect 29043 39080 29055 39083
rect 29086 39080 29092 39092
rect 29043 39052 29092 39080
rect 29043 39049 29055 39052
rect 28997 39043 29055 39049
rect 29086 39040 29092 39052
rect 29144 39040 29150 39092
rect 29822 39040 29828 39092
rect 29880 39080 29886 39092
rect 29880 39052 30696 39080
rect 29880 39040 29886 39052
rect 2406 39012 2412 39024
rect 2367 38984 2412 39012
rect 2406 38972 2412 38984
rect 2464 38972 2470 39024
rect 22830 38972 22836 39024
rect 22888 39012 22894 39024
rect 22888 38984 30420 39012
rect 22888 38972 22894 38984
rect 2222 38944 2228 38956
rect 2183 38916 2228 38944
rect 2222 38904 2228 38916
rect 2280 38904 2286 38956
rect 20901 38947 20959 38953
rect 20901 38913 20913 38947
rect 20947 38913 20959 38947
rect 20901 38907 20959 38913
rect 20993 38947 21051 38953
rect 20993 38913 21005 38947
rect 21039 38913 21051 38947
rect 20993 38907 21051 38913
rect 2774 38876 2780 38888
rect 2735 38848 2780 38876
rect 2774 38836 2780 38848
rect 2832 38836 2838 38888
rect 20916 38808 20944 38907
rect 21008 38876 21036 38907
rect 21082 38904 21088 38956
rect 21140 38944 21146 38956
rect 21269 38947 21327 38953
rect 21140 38916 21185 38944
rect 21140 38904 21146 38916
rect 21269 38913 21281 38947
rect 21315 38913 21327 38947
rect 21269 38907 21327 38913
rect 22005 38947 22063 38953
rect 22005 38913 22017 38947
rect 22051 38944 22063 38947
rect 22094 38944 22100 38956
rect 22051 38916 22100 38944
rect 22051 38913 22063 38916
rect 22005 38907 22063 38913
rect 21174 38876 21180 38888
rect 21008 38848 21180 38876
rect 21174 38836 21180 38848
rect 21232 38836 21238 38888
rect 21284 38876 21312 38907
rect 22094 38904 22100 38916
rect 22152 38904 22158 38956
rect 22370 38944 22376 38956
rect 22204 38916 22376 38944
rect 22204 38876 22232 38916
rect 22370 38904 22376 38916
rect 22428 38904 22434 38956
rect 22646 38904 22652 38956
rect 22704 38944 22710 38956
rect 22741 38947 22799 38953
rect 22741 38944 22753 38947
rect 22704 38916 22753 38944
rect 22704 38904 22710 38916
rect 22741 38913 22753 38916
rect 22787 38913 22799 38947
rect 23382 38944 23388 38956
rect 22741 38907 22799 38913
rect 22848 38916 23388 38944
rect 21284 38848 22232 38876
rect 22278 38836 22284 38888
rect 22336 38876 22342 38888
rect 22848 38876 22876 38916
rect 23382 38904 23388 38916
rect 23440 38904 23446 38956
rect 23842 38944 23848 38956
rect 23803 38916 23848 38944
rect 23842 38904 23848 38916
rect 23900 38904 23906 38956
rect 27614 38904 27620 38956
rect 27672 38944 27678 38956
rect 27985 38947 28043 38953
rect 27985 38944 27997 38947
rect 27672 38916 27997 38944
rect 27672 38904 27678 38916
rect 27985 38913 27997 38916
rect 28031 38913 28043 38947
rect 27985 38907 28043 38913
rect 28261 38947 28319 38953
rect 28261 38913 28273 38947
rect 28307 38944 28319 38947
rect 29457 38947 29515 38953
rect 29457 38944 29469 38947
rect 28307 38916 29469 38944
rect 28307 38913 28319 38916
rect 28261 38907 28319 38913
rect 29457 38913 29469 38916
rect 29503 38913 29515 38947
rect 29457 38907 29515 38913
rect 29546 38904 29552 38956
rect 29604 38944 29610 38956
rect 29641 38947 29699 38953
rect 29641 38944 29653 38947
rect 29604 38916 29653 38944
rect 29604 38904 29610 38916
rect 29641 38913 29653 38916
rect 29687 38913 29699 38947
rect 29641 38907 29699 38913
rect 29917 38947 29975 38953
rect 29917 38913 29929 38947
rect 29963 38944 29975 38947
rect 30006 38944 30012 38956
rect 29963 38916 30012 38944
rect 29963 38913 29975 38916
rect 29917 38907 29975 38913
rect 30006 38904 30012 38916
rect 30064 38904 30070 38956
rect 30101 38947 30159 38953
rect 30101 38913 30113 38947
rect 30147 38944 30159 38947
rect 30190 38944 30196 38956
rect 30147 38916 30196 38944
rect 30147 38913 30159 38916
rect 30101 38907 30159 38913
rect 30190 38904 30196 38916
rect 30248 38904 30254 38956
rect 22336 38848 22876 38876
rect 23017 38879 23075 38885
rect 22336 38836 22342 38848
rect 23017 38845 23029 38879
rect 23063 38876 23075 38879
rect 23063 38848 23520 38876
rect 23063 38845 23075 38848
rect 23017 38839 23075 38845
rect 20990 38808 20996 38820
rect 20916 38780 20996 38808
rect 20990 38768 20996 38780
rect 21048 38768 21054 38820
rect 22833 38811 22891 38817
rect 22833 38777 22845 38811
rect 22879 38808 22891 38811
rect 23198 38808 23204 38820
rect 22879 38780 23204 38808
rect 22879 38777 22891 38780
rect 22833 38771 22891 38777
rect 23198 38768 23204 38780
rect 23256 38768 23262 38820
rect 23492 38808 23520 38848
rect 24394 38836 24400 38888
rect 24452 38876 24458 38888
rect 24581 38879 24639 38885
rect 24581 38876 24593 38879
rect 24452 38848 24593 38876
rect 24452 38836 24458 38848
rect 24581 38845 24593 38848
rect 24627 38845 24639 38879
rect 24581 38839 24639 38845
rect 24670 38836 24676 38888
rect 24728 38876 24734 38888
rect 24857 38879 24915 38885
rect 24857 38876 24869 38879
rect 24728 38848 24869 38876
rect 24728 38836 24734 38848
rect 24857 38845 24869 38848
rect 24903 38845 24915 38879
rect 24857 38839 24915 38845
rect 23842 38808 23848 38820
rect 23492 38780 23848 38808
rect 23842 38768 23848 38780
rect 23900 38808 23906 38820
rect 24688 38808 24716 38836
rect 23900 38780 24716 38808
rect 30392 38808 30420 38984
rect 30466 38972 30472 39024
rect 30524 39012 30530 39024
rect 30561 39015 30619 39021
rect 30561 39012 30573 39015
rect 30524 38984 30573 39012
rect 30524 38972 30530 38984
rect 30561 38981 30573 38984
rect 30607 38981 30619 39015
rect 30668 39012 30696 39052
rect 30742 39040 30748 39092
rect 30800 39089 30806 39092
rect 30800 39083 30819 39089
rect 30807 39080 30819 39083
rect 31018 39080 31024 39092
rect 30807 39052 31024 39080
rect 30807 39049 30819 39052
rect 30800 39043 30819 39049
rect 30800 39040 30806 39043
rect 31018 39040 31024 39052
rect 31076 39040 31082 39092
rect 31478 39080 31484 39092
rect 31439 39052 31484 39080
rect 31478 39040 31484 39052
rect 31536 39040 31542 39092
rect 33042 39080 33048 39092
rect 33003 39052 33048 39080
rect 33042 39040 33048 39052
rect 33100 39040 33106 39092
rect 34333 39083 34391 39089
rect 34333 39049 34345 39083
rect 34379 39080 34391 39083
rect 35434 39080 35440 39092
rect 34379 39052 35440 39080
rect 34379 39049 34391 39052
rect 34333 39043 34391 39049
rect 35434 39040 35440 39052
rect 35492 39040 35498 39092
rect 37642 39080 37648 39092
rect 37476 39052 37648 39080
rect 30668 38984 31616 39012
rect 30561 38975 30619 38981
rect 30834 38904 30840 38956
rect 30892 38944 30898 38956
rect 31588 38953 31616 38984
rect 31754 38972 31760 39024
rect 31812 39012 31818 39024
rect 32306 39012 32312 39024
rect 31812 38984 32312 39012
rect 31812 38972 31818 38984
rect 32306 38972 32312 38984
rect 32364 39012 32370 39024
rect 32674 39012 32680 39024
rect 32364 38984 32444 39012
rect 32635 38984 32680 39012
rect 32364 38972 32370 38984
rect 32416 38953 32444 38984
rect 32674 38972 32680 38984
rect 32732 38972 32738 39024
rect 32769 39015 32827 39021
rect 32769 38981 32781 39015
rect 32815 39012 32827 39015
rect 36078 39012 36084 39024
rect 32815 38984 36084 39012
rect 32815 38981 32827 38984
rect 32769 38975 32827 38981
rect 36078 38972 36084 38984
rect 36136 38972 36142 39024
rect 31389 38950 31447 38953
rect 31328 38947 31447 38950
rect 31328 38944 31401 38947
rect 30892 38922 31401 38944
rect 30892 38916 31356 38922
rect 30892 38904 30898 38916
rect 31389 38913 31401 38922
rect 31435 38913 31447 38947
rect 31389 38907 31447 38913
rect 31573 38947 31631 38953
rect 31573 38913 31585 38947
rect 31619 38944 31631 38947
rect 32401 38947 32459 38953
rect 31619 38916 32352 38944
rect 31619 38913 31631 38916
rect 31573 38907 31631 38913
rect 32324 38876 32352 38916
rect 32401 38913 32413 38947
rect 32447 38913 32459 38947
rect 32401 38907 32459 38913
rect 32490 38904 32496 38956
rect 32548 38944 32554 38956
rect 32907 38947 32965 38953
rect 32548 38916 32593 38944
rect 32548 38904 32554 38916
rect 32907 38913 32919 38947
rect 32953 38944 32965 38947
rect 33318 38944 33324 38956
rect 32953 38916 33324 38944
rect 32953 38913 32965 38916
rect 32907 38907 32965 38913
rect 33318 38904 33324 38916
rect 33376 38904 33382 38956
rect 33505 38947 33563 38953
rect 33505 38913 33517 38947
rect 33551 38913 33563 38947
rect 33505 38907 33563 38913
rect 33520 38876 33548 38907
rect 33778 38904 33784 38956
rect 33836 38944 33842 38956
rect 34517 38947 34575 38953
rect 34517 38944 34529 38947
rect 33836 38916 34529 38944
rect 33836 38904 33842 38916
rect 34517 38913 34529 38916
rect 34563 38944 34575 38947
rect 34882 38944 34888 38956
rect 34563 38916 34888 38944
rect 34563 38913 34575 38916
rect 34517 38907 34575 38913
rect 34882 38904 34888 38916
rect 34940 38904 34946 38956
rect 35345 38947 35403 38953
rect 35345 38913 35357 38947
rect 35391 38913 35403 38947
rect 35345 38907 35403 38913
rect 35529 38947 35587 38953
rect 35529 38913 35541 38947
rect 35575 38944 35587 38947
rect 37274 38944 37280 38956
rect 35575 38916 37136 38944
rect 37235 38916 37280 38944
rect 35575 38913 35587 38916
rect 35529 38907 35587 38913
rect 32324 38848 33548 38876
rect 34146 38836 34152 38888
rect 34204 38876 34210 38888
rect 34609 38879 34667 38885
rect 34609 38876 34621 38879
rect 34204 38848 34621 38876
rect 34204 38836 34210 38848
rect 34609 38845 34621 38848
rect 34655 38845 34667 38879
rect 34609 38839 34667 38845
rect 34701 38879 34759 38885
rect 34701 38845 34713 38879
rect 34747 38845 34759 38879
rect 34701 38839 34759 38845
rect 34793 38879 34851 38885
rect 34793 38845 34805 38879
rect 34839 38845 34851 38879
rect 35360 38876 35388 38907
rect 35710 38876 35716 38888
rect 35360 38848 35716 38876
rect 34793 38839 34851 38845
rect 32490 38808 32496 38820
rect 30392 38780 32496 38808
rect 23900 38768 23906 38780
rect 32490 38768 32496 38780
rect 32548 38768 32554 38820
rect 33594 38808 33600 38820
rect 33555 38780 33600 38808
rect 33594 38768 33600 38780
rect 33652 38768 33658 38820
rect 34238 38768 34244 38820
rect 34296 38808 34302 38820
rect 34716 38808 34744 38839
rect 34296 38780 34744 38808
rect 34296 38768 34302 38780
rect 19518 38700 19524 38752
rect 19576 38740 19582 38752
rect 20625 38743 20683 38749
rect 20625 38740 20637 38743
rect 19576 38712 20637 38740
rect 19576 38700 19582 38712
rect 20625 38709 20637 38712
rect 20671 38709 20683 38743
rect 20625 38703 20683 38709
rect 20806 38700 20812 38752
rect 20864 38740 20870 38752
rect 21821 38743 21879 38749
rect 21821 38740 21833 38743
rect 20864 38712 21833 38740
rect 20864 38700 20870 38712
rect 21821 38709 21833 38712
rect 21867 38709 21879 38743
rect 22186 38740 22192 38752
rect 22147 38712 22192 38740
rect 21821 38703 21879 38709
rect 22186 38700 22192 38712
rect 22244 38700 22250 38752
rect 22922 38700 22928 38752
rect 22980 38740 22986 38752
rect 23934 38740 23940 38752
rect 22980 38712 23025 38740
rect 23895 38712 23940 38740
rect 22980 38700 22986 38712
rect 23934 38700 23940 38712
rect 23992 38700 23998 38752
rect 30006 38700 30012 38752
rect 30064 38740 30070 38752
rect 30745 38743 30803 38749
rect 30745 38740 30757 38743
rect 30064 38712 30757 38740
rect 30064 38700 30070 38712
rect 30745 38709 30757 38712
rect 30791 38709 30803 38743
rect 30926 38740 30932 38752
rect 30887 38712 30932 38740
rect 30745 38703 30803 38709
rect 30926 38700 30932 38712
rect 30984 38700 30990 38752
rect 32508 38740 32536 38768
rect 34808 38752 34836 38839
rect 35710 38836 35716 38848
rect 35768 38836 35774 38888
rect 37108 38876 37136 38916
rect 37274 38904 37280 38916
rect 37332 38904 37338 38956
rect 37476 38953 37504 39052
rect 37642 39040 37648 39052
rect 37700 39040 37706 39092
rect 38470 39040 38476 39092
rect 38528 39080 38534 39092
rect 40218 39080 40224 39092
rect 38528 39052 40224 39080
rect 38528 39040 38534 39052
rect 40218 39040 40224 39052
rect 40276 39080 40282 39092
rect 40276 39052 40366 39080
rect 40276 39040 40282 39052
rect 40494 39040 40500 39092
rect 40552 39080 40558 39092
rect 40957 39083 41015 39089
rect 40957 39080 40969 39083
rect 40552 39052 40969 39080
rect 40552 39040 40558 39052
rect 40957 39049 40969 39052
rect 41003 39049 41015 39083
rect 40957 39043 41015 39049
rect 43441 39083 43499 39089
rect 43441 39049 43453 39083
rect 43487 39080 43499 39083
rect 45646 39080 45652 39092
rect 43487 39052 45652 39080
rect 43487 39049 43499 39052
rect 43441 39043 43499 39049
rect 45646 39040 45652 39052
rect 45704 39040 45710 39092
rect 46014 39040 46020 39092
rect 46072 39040 46078 39092
rect 49234 39040 49240 39092
rect 49292 39080 49298 39092
rect 50157 39083 50215 39089
rect 50157 39080 50169 39083
rect 49292 39052 50169 39080
rect 49292 39040 49298 39052
rect 50157 39049 50169 39052
rect 50203 39080 50215 39083
rect 50939 39083 50997 39089
rect 50939 39080 50951 39083
rect 50203 39052 50951 39080
rect 50203 39049 50215 39052
rect 50157 39043 50215 39049
rect 50939 39049 50951 39052
rect 50985 39049 50997 39083
rect 52086 39080 52092 39092
rect 52047 39052 52092 39080
rect 50939 39043 50997 39049
rect 52086 39040 52092 39052
rect 52144 39040 52150 39092
rect 53466 39080 53472 39092
rect 53427 39052 53472 39080
rect 53466 39040 53472 39052
rect 53524 39040 53530 39092
rect 37553 39015 37611 39021
rect 37553 38981 37565 39015
rect 37599 39012 37611 39015
rect 39390 39012 39396 39024
rect 37599 38984 39396 39012
rect 37599 38981 37611 38984
rect 37553 38975 37611 38981
rect 39390 38972 39396 38984
rect 39448 38972 39454 39024
rect 37461 38947 37519 38953
rect 37461 38913 37473 38947
rect 37507 38913 37519 38947
rect 37461 38907 37519 38913
rect 37645 38947 37703 38953
rect 37645 38913 37657 38947
rect 37691 38944 37703 38947
rect 37826 38944 37832 38956
rect 37691 38916 37832 38944
rect 37691 38913 37703 38916
rect 37645 38907 37703 38913
rect 37826 38904 37832 38916
rect 37884 38904 37890 38956
rect 38378 38944 38384 38956
rect 38339 38916 38384 38944
rect 38378 38904 38384 38916
rect 38436 38904 38442 38956
rect 38562 38944 38568 38956
rect 38523 38916 38568 38944
rect 38562 38904 38568 38916
rect 38620 38904 38626 38956
rect 39764 38947 39822 38953
rect 39592 38944 39712 38947
rect 39592 38942 39728 38944
rect 39764 38942 39776 38947
rect 39592 38919 39776 38942
rect 39482 38876 39488 38888
rect 37108 38848 39488 38876
rect 39482 38836 39488 38848
rect 39540 38876 39546 38888
rect 39592 38876 39620 38919
rect 39684 38916 39776 38919
rect 39700 38914 39776 38916
rect 39764 38913 39776 38914
rect 39810 38913 39822 38947
rect 39764 38907 39822 38913
rect 39853 38947 39911 38953
rect 39853 38913 39865 38947
rect 39899 38913 39911 38947
rect 40034 38944 40040 38956
rect 39995 38916 40040 38944
rect 39853 38907 39911 38913
rect 39868 38876 39896 38907
rect 40034 38904 40040 38916
rect 40092 38904 40098 38956
rect 40139 38947 40197 38953
rect 40139 38913 40151 38947
rect 40185 38944 40197 38947
rect 40233 38944 40261 39040
rect 41598 38972 41604 39024
rect 41656 39012 41662 39024
rect 41693 39015 41751 39021
rect 41693 39012 41705 39015
rect 41656 38984 41705 39012
rect 41656 38972 41662 38984
rect 41693 38981 41705 38984
rect 41739 39012 41751 39015
rect 42150 39012 42156 39024
rect 41739 38984 42156 39012
rect 41739 38981 41751 38984
rect 41693 38975 41751 38981
rect 42150 38972 42156 38984
rect 42208 38972 42214 39024
rect 45370 39012 45376 39024
rect 43548 38984 43852 39012
rect 40586 38944 40592 38956
rect 40185 38916 40261 38944
rect 40499 38916 40592 38944
rect 40185 38913 40197 38916
rect 40139 38907 40197 38913
rect 40586 38904 40592 38916
rect 40644 38944 40650 38956
rect 40644 38916 41460 38944
rect 40644 38904 40650 38916
rect 39540 38848 39620 38876
rect 39684 38848 39896 38876
rect 40681 38879 40739 38885
rect 39540 38836 39546 38848
rect 39684 38820 39712 38848
rect 40681 38845 40693 38879
rect 40727 38845 40739 38879
rect 41432 38876 41460 38916
rect 41506 38904 41512 38956
rect 41564 38944 41570 38956
rect 43548 38944 43576 38984
rect 41564 38916 43576 38944
rect 43625 38947 43683 38953
rect 41564 38904 41570 38916
rect 43625 38913 43637 38947
rect 43671 38913 43683 38947
rect 43625 38907 43683 38913
rect 43717 38947 43775 38953
rect 43717 38913 43729 38947
rect 43763 38913 43775 38947
rect 43717 38907 43775 38913
rect 43530 38876 43536 38888
rect 41432 38848 43536 38876
rect 40681 38839 40739 38845
rect 35618 38768 35624 38820
rect 35676 38808 35682 38820
rect 39022 38808 39028 38820
rect 35676 38780 39028 38808
rect 35676 38768 35682 38780
rect 39022 38768 39028 38780
rect 39080 38768 39086 38820
rect 39390 38768 39396 38820
rect 39448 38808 39454 38820
rect 39577 38811 39635 38817
rect 39577 38808 39589 38811
rect 39448 38780 39589 38808
rect 39448 38768 39454 38780
rect 39577 38777 39589 38780
rect 39623 38777 39635 38811
rect 39577 38771 39635 38777
rect 39666 38768 39672 38820
rect 39724 38768 39730 38820
rect 40126 38768 40132 38820
rect 40184 38808 40190 38820
rect 40696 38808 40724 38839
rect 43530 38836 43536 38848
rect 43588 38836 43594 38888
rect 40184 38780 40724 38808
rect 40184 38768 40190 38780
rect 34330 38740 34336 38752
rect 32508 38712 34336 38740
rect 34330 38700 34336 38712
rect 34388 38700 34394 38752
rect 34790 38700 34796 38752
rect 34848 38700 34854 38752
rect 35345 38743 35403 38749
rect 35345 38709 35357 38743
rect 35391 38740 35403 38743
rect 35526 38740 35532 38752
rect 35391 38712 35532 38740
rect 35391 38709 35403 38712
rect 35345 38703 35403 38709
rect 35526 38700 35532 38712
rect 35584 38700 35590 38752
rect 37642 38700 37648 38752
rect 37700 38740 37706 38752
rect 37829 38743 37887 38749
rect 37829 38740 37841 38743
rect 37700 38712 37841 38740
rect 37700 38700 37706 38712
rect 37829 38709 37841 38712
rect 37875 38709 37887 38743
rect 40586 38740 40592 38752
rect 40547 38712 40592 38740
rect 37829 38703 37887 38709
rect 40586 38700 40592 38712
rect 40644 38700 40650 38752
rect 43640 38740 43668 38907
rect 43732 38808 43760 38907
rect 43824 38876 43852 38984
rect 43916 38984 45376 39012
rect 43916 38953 43944 38984
rect 45370 38972 45376 38984
rect 45428 38972 45434 39024
rect 43901 38947 43959 38953
rect 43901 38913 43913 38947
rect 43947 38913 43959 38947
rect 43901 38907 43959 38913
rect 43993 38947 44051 38953
rect 43993 38913 44005 38947
rect 44039 38944 44051 38947
rect 44358 38944 44364 38956
rect 44039 38916 44364 38944
rect 44039 38913 44051 38916
rect 43993 38907 44051 38913
rect 44008 38876 44036 38907
rect 44358 38904 44364 38916
rect 44416 38904 44422 38956
rect 44726 38944 44732 38956
rect 44687 38916 44732 38944
rect 44726 38904 44732 38916
rect 44784 38904 44790 38956
rect 45002 38944 45008 38956
rect 44963 38916 45008 38944
rect 45002 38904 45008 38916
rect 45060 38904 45066 38956
rect 45189 38947 45247 38953
rect 45189 38913 45201 38947
rect 45235 38944 45247 38947
rect 45462 38944 45468 38956
rect 45235 38916 45468 38944
rect 45235 38913 45247 38916
rect 45189 38907 45247 38913
rect 43824 38848 44036 38876
rect 44082 38836 44088 38888
rect 44140 38876 44146 38888
rect 45204 38876 45232 38907
rect 45462 38904 45468 38916
rect 45520 38904 45526 38956
rect 45830 38904 45836 38956
rect 45888 38944 45894 38956
rect 46032 38953 46060 39040
rect 48498 39012 48504 39024
rect 48411 38984 48504 39012
rect 48498 38972 48504 38984
rect 48556 39012 48562 39024
rect 48774 39012 48780 39024
rect 48556 38984 48780 39012
rect 48556 38972 48562 38984
rect 48774 38972 48780 38984
rect 48832 38972 48838 39024
rect 49973 39015 50031 39021
rect 49973 38981 49985 39015
rect 50019 39012 50031 39015
rect 50019 38984 51074 39012
rect 50019 38981 50031 38984
rect 49973 38975 50031 38981
rect 45925 38947 45983 38953
rect 45925 38944 45937 38947
rect 45888 38916 45937 38944
rect 45888 38904 45894 38916
rect 45925 38913 45937 38916
rect 45971 38913 45983 38947
rect 45925 38907 45983 38913
rect 46017 38947 46075 38953
rect 46017 38913 46029 38947
rect 46063 38913 46075 38947
rect 46017 38907 46075 38913
rect 46109 38947 46167 38953
rect 46109 38913 46121 38947
rect 46155 38913 46167 38947
rect 46109 38907 46167 38913
rect 46293 38947 46351 38953
rect 46293 38913 46305 38947
rect 46339 38944 46351 38947
rect 46845 38947 46903 38953
rect 46339 38916 46428 38944
rect 46339 38913 46351 38916
rect 46293 38907 46351 38913
rect 44140 38848 45232 38876
rect 44140 38836 44146 38848
rect 45554 38836 45560 38888
rect 45612 38876 45618 38888
rect 46124 38876 46152 38907
rect 45612 38848 46152 38876
rect 46400 38876 46428 38916
rect 46845 38913 46857 38947
rect 46891 38944 46903 38947
rect 48038 38944 48044 38956
rect 46891 38916 48044 38944
rect 46891 38913 46903 38916
rect 46845 38907 46903 38913
rect 48038 38904 48044 38916
rect 48096 38904 48102 38956
rect 48317 38947 48375 38953
rect 48317 38913 48329 38947
rect 48363 38913 48375 38947
rect 48317 38907 48375 38913
rect 49329 38947 49387 38953
rect 49329 38913 49341 38947
rect 49375 38944 49387 38947
rect 50249 38947 50307 38953
rect 49375 38916 50200 38944
rect 49375 38913 49387 38916
rect 49329 38907 49387 38913
rect 46934 38876 46940 38888
rect 46400 38848 46940 38876
rect 45612 38836 45618 38848
rect 44726 38808 44732 38820
rect 43732 38780 44732 38808
rect 44726 38768 44732 38780
rect 44784 38768 44790 38820
rect 44821 38811 44879 38817
rect 44821 38777 44833 38811
rect 44867 38808 44879 38811
rect 46290 38808 46296 38820
rect 44867 38780 46296 38808
rect 44867 38777 44879 38780
rect 44821 38771 44879 38777
rect 46290 38768 46296 38780
rect 46348 38768 46354 38820
rect 44266 38740 44272 38752
rect 43640 38712 44272 38740
rect 44266 38700 44272 38712
rect 44324 38700 44330 38752
rect 44450 38740 44456 38752
rect 44411 38712 44456 38740
rect 44450 38700 44456 38712
rect 44508 38700 44514 38752
rect 44634 38700 44640 38752
rect 44692 38740 44698 38752
rect 44913 38743 44971 38749
rect 44913 38740 44925 38743
rect 44692 38712 44925 38740
rect 44692 38700 44698 38712
rect 44913 38709 44925 38712
rect 44959 38740 44971 38743
rect 45649 38743 45707 38749
rect 45649 38740 45661 38743
rect 44959 38712 45661 38740
rect 44959 38709 44971 38712
rect 44913 38703 44971 38709
rect 45649 38709 45661 38712
rect 45695 38709 45707 38743
rect 45649 38703 45707 38709
rect 45738 38700 45744 38752
rect 45796 38740 45802 38752
rect 46400 38740 46428 38848
rect 46934 38836 46940 38848
rect 46992 38836 46998 38888
rect 48332 38808 48360 38907
rect 48406 38836 48412 38888
rect 48464 38876 48470 38888
rect 48958 38876 48964 38888
rect 48464 38848 48964 38876
rect 48464 38836 48470 38848
rect 48958 38836 48964 38848
rect 49016 38876 49022 38888
rect 49421 38879 49479 38885
rect 49421 38876 49433 38879
rect 49016 38848 49433 38876
rect 49016 38836 49022 38848
rect 49421 38845 49433 38848
rect 49467 38845 49479 38879
rect 49421 38839 49479 38845
rect 49694 38836 49700 38888
rect 49752 38876 49758 38888
rect 49878 38876 49884 38888
rect 49752 38848 49884 38876
rect 49752 38836 49758 38848
rect 49878 38836 49884 38848
rect 49936 38836 49942 38888
rect 50172 38876 50200 38916
rect 50249 38913 50261 38947
rect 50295 38944 50307 38947
rect 50614 38944 50620 38956
rect 50295 38916 50620 38944
rect 50295 38913 50307 38916
rect 50249 38907 50307 38913
rect 50614 38904 50620 38916
rect 50672 38904 50678 38956
rect 50706 38876 50712 38888
rect 50172 38848 50712 38876
rect 50706 38836 50712 38848
rect 50764 38836 50770 38888
rect 51046 38876 51074 38984
rect 51997 38947 52055 38953
rect 51997 38913 52009 38947
rect 52043 38913 52055 38947
rect 52178 38944 52184 38956
rect 52139 38916 52184 38944
rect 51997 38907 52055 38913
rect 51902 38876 51908 38888
rect 51046 38848 51908 38876
rect 51902 38836 51908 38848
rect 51960 38836 51966 38888
rect 49973 38811 50031 38817
rect 48332 38780 49740 38808
rect 46934 38740 46940 38752
rect 45796 38712 46428 38740
rect 46895 38712 46940 38740
rect 45796 38700 45802 38712
rect 46934 38700 46940 38712
rect 46992 38700 46998 38752
rect 48682 38700 48688 38752
rect 48740 38740 48746 38752
rect 48958 38740 48964 38752
rect 48740 38712 48964 38740
rect 48740 38700 48746 38712
rect 48958 38700 48964 38712
rect 49016 38700 49022 38752
rect 49712 38740 49740 38780
rect 49973 38777 49985 38811
rect 50019 38808 50031 38811
rect 52012 38808 52040 38907
rect 52178 38904 52184 38916
rect 52236 38904 52242 38956
rect 53282 38944 53288 38956
rect 53243 38916 53288 38944
rect 53282 38904 53288 38916
rect 53340 38904 53346 38956
rect 53101 38879 53159 38885
rect 53101 38845 53113 38879
rect 53147 38876 53159 38879
rect 53650 38876 53656 38888
rect 53147 38848 53656 38876
rect 53147 38845 53159 38848
rect 53101 38839 53159 38845
rect 53650 38836 53656 38848
rect 53708 38836 53714 38888
rect 50019 38780 52040 38808
rect 50019 38777 50031 38780
rect 49973 38771 50031 38777
rect 51442 38740 51448 38752
rect 49712 38712 51448 38740
rect 51442 38700 51448 38712
rect 51500 38740 51506 38752
rect 51718 38740 51724 38752
rect 51500 38712 51724 38740
rect 51500 38700 51506 38712
rect 51718 38700 51724 38712
rect 51776 38700 51782 38752
rect 56594 38700 56600 38752
rect 56652 38740 56658 38752
rect 58069 38743 58127 38749
rect 58069 38740 58081 38743
rect 56652 38712 58081 38740
rect 56652 38700 56658 38712
rect 58069 38709 58081 38712
rect 58115 38709 58127 38743
rect 58069 38703 58127 38709
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 21174 38496 21180 38548
rect 21232 38536 21238 38548
rect 23934 38536 23940 38548
rect 21232 38508 23940 38536
rect 21232 38496 21238 38508
rect 19245 38335 19303 38341
rect 19245 38301 19257 38335
rect 19291 38332 19303 38335
rect 20622 38332 20628 38344
rect 19291 38304 20628 38332
rect 19291 38301 19303 38304
rect 19245 38295 19303 38301
rect 20622 38292 20628 38304
rect 20680 38292 20686 38344
rect 19518 38273 19524 38276
rect 19512 38264 19524 38273
rect 19479 38236 19524 38264
rect 19512 38227 19524 38236
rect 19518 38224 19524 38227
rect 19576 38224 19582 38276
rect 21744 38264 21772 38508
rect 23934 38496 23940 38508
rect 23992 38496 23998 38548
rect 29362 38496 29368 38548
rect 29420 38536 29426 38548
rect 29549 38539 29607 38545
rect 29549 38536 29561 38539
rect 29420 38508 29561 38536
rect 29420 38496 29426 38508
rect 29549 38505 29561 38508
rect 29595 38505 29607 38539
rect 29549 38499 29607 38505
rect 29656 38508 34744 38536
rect 22278 38468 22284 38480
rect 21908 38440 22284 38468
rect 21908 38341 21936 38440
rect 22278 38428 22284 38440
rect 22336 38428 22342 38480
rect 24394 38428 24400 38480
rect 24452 38468 24458 38480
rect 26694 38468 26700 38480
rect 24452 38440 24992 38468
rect 26607 38440 26700 38468
rect 24452 38428 24458 38440
rect 22741 38403 22799 38409
rect 22741 38400 22753 38403
rect 22204 38372 22753 38400
rect 21908 38335 21971 38341
rect 21908 38301 21925 38335
rect 21959 38301 21971 38335
rect 22005 38335 22063 38341
rect 22005 38310 22017 38335
rect 21913 38295 21971 38301
rect 22001 38301 22017 38310
rect 22051 38301 22063 38335
rect 22001 38295 22063 38301
rect 22118 38332 22176 38338
rect 22118 38298 22130 38332
rect 22164 38329 22176 38332
rect 22204 38329 22232 38372
rect 22741 38369 22753 38372
rect 22787 38369 22799 38403
rect 22741 38363 22799 38369
rect 24578 38360 24584 38412
rect 24636 38400 24642 38412
rect 24964 38409 24992 38440
rect 26694 38428 26700 38440
rect 26752 38468 26758 38480
rect 27522 38468 27528 38480
rect 26752 38440 27528 38468
rect 26752 38428 26758 38440
rect 27522 38428 27528 38440
rect 27580 38428 27586 38480
rect 27706 38428 27712 38480
rect 27764 38468 27770 38480
rect 29656 38468 29684 38508
rect 27764 38440 29684 38468
rect 27764 38428 27770 38440
rect 30282 38428 30288 38480
rect 30340 38468 30346 38480
rect 34716 38468 34744 38508
rect 34790 38496 34796 38548
rect 34848 38536 34854 38548
rect 35713 38539 35771 38545
rect 35713 38536 35725 38539
rect 34848 38508 35725 38536
rect 34848 38496 34854 38508
rect 35713 38505 35725 38508
rect 35759 38505 35771 38539
rect 35713 38499 35771 38505
rect 36722 38496 36728 38548
rect 36780 38536 36786 38548
rect 38473 38539 38531 38545
rect 36780 38508 38424 38536
rect 36780 38496 36786 38508
rect 37550 38468 37556 38480
rect 30340 38440 33916 38468
rect 34716 38440 35296 38468
rect 30340 38428 30346 38440
rect 24857 38403 24915 38409
rect 24857 38400 24869 38403
rect 24636 38372 24869 38400
rect 24636 38360 24642 38372
rect 24857 38369 24869 38372
rect 24903 38369 24915 38403
rect 24857 38363 24915 38369
rect 24949 38403 25007 38409
rect 24949 38369 24961 38403
rect 24995 38369 25007 38403
rect 30926 38400 30932 38412
rect 24949 38363 25007 38369
rect 30024 38372 30932 38400
rect 22164 38301 22232 38329
rect 22281 38335 22339 38341
rect 22281 38301 22293 38335
rect 22327 38332 22339 38335
rect 22370 38332 22376 38344
rect 22327 38304 22376 38332
rect 22327 38301 22339 38304
rect 22164 38298 22176 38301
rect 22001 38282 22048 38295
rect 22118 38292 22176 38298
rect 22281 38295 22339 38301
rect 22370 38292 22376 38304
rect 22428 38292 22434 38344
rect 22646 38292 22652 38344
rect 22704 38292 22710 38344
rect 22922 38332 22928 38344
rect 22883 38304 22928 38332
rect 22922 38292 22928 38304
rect 22980 38292 22986 38344
rect 23198 38332 23204 38344
rect 23159 38304 23204 38332
rect 23198 38292 23204 38304
rect 23256 38292 23262 38344
rect 24486 38292 24492 38344
rect 24544 38332 24550 38344
rect 24765 38335 24823 38341
rect 24765 38332 24777 38335
rect 24544 38304 24777 38332
rect 24544 38292 24550 38304
rect 24765 38301 24777 38304
rect 24811 38301 24823 38335
rect 25038 38332 25044 38344
rect 24999 38304 25044 38332
rect 24765 38295 24823 38301
rect 25038 38292 25044 38304
rect 25096 38292 25102 38344
rect 28534 38292 28540 38344
rect 28592 38332 28598 38344
rect 30024 38341 30052 38372
rect 30926 38360 30932 38372
rect 30984 38360 30990 38412
rect 31110 38360 31116 38412
rect 31168 38400 31174 38412
rect 32401 38403 32459 38409
rect 32401 38400 32413 38403
rect 31168 38372 32413 38400
rect 31168 38360 31174 38372
rect 32401 38369 32413 38372
rect 32447 38369 32459 38403
rect 32401 38363 32459 38369
rect 29733 38335 29791 38341
rect 29733 38332 29745 38335
rect 28592 38304 29745 38332
rect 28592 38292 28598 38304
rect 29733 38301 29745 38304
rect 29779 38301 29791 38335
rect 29733 38295 29791 38301
rect 30009 38335 30067 38341
rect 30009 38301 30021 38335
rect 30055 38301 30067 38335
rect 30009 38295 30067 38301
rect 30193 38335 30251 38341
rect 30193 38301 30205 38335
rect 30239 38332 30251 38335
rect 30374 38332 30380 38344
rect 30239 38304 30380 38332
rect 30239 38301 30251 38304
rect 30193 38295 30251 38301
rect 22001 38264 22029 38282
rect 21744 38236 22029 38264
rect 22462 38224 22468 38276
rect 22520 38264 22526 38276
rect 22664 38264 22692 38292
rect 23109 38267 23167 38273
rect 23109 38264 23121 38267
rect 22520 38236 23121 38264
rect 22520 38224 22526 38236
rect 23109 38233 23121 38236
rect 23155 38233 23167 38267
rect 26510 38264 26516 38276
rect 26471 38236 26516 38264
rect 23109 38227 23167 38233
rect 26510 38224 26516 38236
rect 26568 38224 26574 38276
rect 29748 38264 29776 38295
rect 30374 38292 30380 38304
rect 30432 38292 30438 38344
rect 30466 38292 30472 38344
rect 30524 38332 30530 38344
rect 30653 38335 30711 38341
rect 30653 38332 30665 38335
rect 30524 38304 30665 38332
rect 30524 38292 30530 38304
rect 30653 38301 30665 38304
rect 30699 38301 30711 38335
rect 30653 38295 30711 38301
rect 30742 38292 30748 38344
rect 30800 38332 30806 38344
rect 31021 38335 31079 38341
rect 31021 38332 31033 38335
rect 30800 38304 31033 38332
rect 30800 38292 30806 38304
rect 31021 38301 31033 38304
rect 31067 38332 31079 38335
rect 32677 38335 32735 38341
rect 31067 38304 31754 38332
rect 31067 38301 31079 38304
rect 31021 38295 31079 38301
rect 30098 38264 30104 38276
rect 29748 38236 30104 38264
rect 30098 38224 30104 38236
rect 30156 38224 30162 38276
rect 30837 38267 30895 38273
rect 30837 38264 30849 38267
rect 30484 38236 30849 38264
rect 20625 38199 20683 38205
rect 20625 38165 20637 38199
rect 20671 38196 20683 38199
rect 20714 38196 20720 38208
rect 20671 38168 20720 38196
rect 20671 38165 20683 38168
rect 20625 38159 20683 38165
rect 20714 38156 20720 38168
rect 20772 38156 20778 38208
rect 21634 38196 21640 38208
rect 21595 38168 21640 38196
rect 21634 38156 21640 38168
rect 21692 38156 21698 38208
rect 22094 38156 22100 38208
rect 22152 38196 22158 38208
rect 22646 38196 22652 38208
rect 22152 38168 22652 38196
rect 22152 38156 22158 38168
rect 22646 38156 22652 38168
rect 22704 38156 22710 38208
rect 24581 38199 24639 38205
rect 24581 38165 24593 38199
rect 24627 38196 24639 38199
rect 25498 38196 25504 38208
rect 24627 38168 25504 38196
rect 24627 38165 24639 38168
rect 24581 38159 24639 38165
rect 25498 38156 25504 38168
rect 25556 38156 25562 38208
rect 29822 38156 29828 38208
rect 29880 38196 29886 38208
rect 30484 38196 30512 38236
rect 30837 38233 30849 38236
rect 30883 38233 30895 38267
rect 30837 38227 30895 38233
rect 31478 38224 31484 38276
rect 31536 38264 31542 38276
rect 31573 38267 31631 38273
rect 31573 38264 31585 38267
rect 31536 38236 31585 38264
rect 31536 38224 31542 38236
rect 31573 38233 31585 38236
rect 31619 38233 31631 38267
rect 31726 38264 31754 38304
rect 32677 38301 32689 38335
rect 32723 38332 32735 38335
rect 33318 38332 33324 38344
rect 32723 38304 33324 38332
rect 32723 38301 32735 38304
rect 32677 38295 32735 38301
rect 33318 38292 33324 38304
rect 33376 38292 33382 38344
rect 33888 38341 33916 38440
rect 34977 38403 35035 38409
rect 34977 38400 34989 38403
rect 34808 38372 34989 38400
rect 33689 38335 33747 38341
rect 33689 38301 33701 38335
rect 33735 38301 33747 38335
rect 33689 38295 33747 38301
rect 33873 38335 33931 38341
rect 33873 38301 33885 38335
rect 33919 38301 33931 38335
rect 33873 38295 33931 38301
rect 33704 38264 33732 38295
rect 34146 38292 34152 38344
rect 34204 38332 34210 38344
rect 34808 38332 34836 38372
rect 34977 38369 34989 38372
rect 35023 38369 35035 38403
rect 35158 38400 35164 38412
rect 35119 38372 35164 38400
rect 34977 38363 35035 38369
rect 35158 38360 35164 38372
rect 35216 38360 35222 38412
rect 35268 38400 35296 38440
rect 36648 38440 37556 38468
rect 36538 38400 36544 38412
rect 35268 38372 36544 38400
rect 34204 38304 34836 38332
rect 34885 38335 34943 38341
rect 34204 38292 34210 38304
rect 34885 38301 34897 38335
rect 34931 38301 34943 38335
rect 34885 38295 34943 38301
rect 35069 38335 35127 38341
rect 35069 38301 35081 38335
rect 35115 38332 35127 38335
rect 35268 38332 35296 38372
rect 35115 38304 35296 38332
rect 35115 38301 35127 38304
rect 35069 38295 35127 38301
rect 31726 38236 33732 38264
rect 33781 38267 33839 38273
rect 31573 38227 31631 38233
rect 33781 38233 33793 38267
rect 33827 38233 33839 38267
rect 33781 38227 33839 38233
rect 29880 38168 30512 38196
rect 29880 38156 29886 38168
rect 31294 38156 31300 38208
rect 31352 38196 31358 38208
rect 31665 38199 31723 38205
rect 31665 38196 31677 38199
rect 31352 38168 31677 38196
rect 31352 38156 31358 38168
rect 31665 38165 31677 38168
rect 31711 38165 31723 38199
rect 33796 38196 33824 38227
rect 34330 38196 34336 38208
rect 33796 38168 34336 38196
rect 31665 38159 31723 38165
rect 34330 38156 34336 38168
rect 34388 38156 34394 38208
rect 34606 38156 34612 38208
rect 34664 38196 34670 38208
rect 34701 38199 34759 38205
rect 34701 38196 34713 38199
rect 34664 38168 34713 38196
rect 34664 38156 34670 38168
rect 34701 38165 34713 38168
rect 34747 38165 34759 38199
rect 34701 38159 34759 38165
rect 34790 38156 34796 38208
rect 34848 38196 34854 38208
rect 34900 38196 34928 38295
rect 35618 38292 35624 38344
rect 35676 38332 35682 38344
rect 35713 38335 35771 38341
rect 35713 38332 35725 38335
rect 35676 38304 35725 38332
rect 35676 38292 35682 38304
rect 35713 38301 35725 38304
rect 35759 38301 35771 38335
rect 35713 38295 35771 38301
rect 35897 38335 35955 38341
rect 35897 38301 35909 38335
rect 35943 38332 35955 38335
rect 36262 38332 36268 38344
rect 35943 38304 36268 38332
rect 35943 38301 35955 38304
rect 35897 38295 35955 38301
rect 36262 38292 36268 38304
rect 36320 38292 36326 38344
rect 36464 38341 36492 38372
rect 36538 38360 36544 38372
rect 36596 38360 36602 38412
rect 36648 38344 36676 38440
rect 37550 38428 37556 38440
rect 37608 38428 37614 38480
rect 38396 38468 38424 38508
rect 38473 38505 38485 38539
rect 38519 38536 38531 38539
rect 38654 38536 38660 38548
rect 38519 38508 38660 38536
rect 38519 38505 38531 38508
rect 38473 38499 38531 38505
rect 38654 38496 38660 38508
rect 38712 38496 38718 38548
rect 41322 38496 41328 38548
rect 41380 38536 41386 38548
rect 41380 38496 41414 38536
rect 44726 38496 44732 38548
rect 44784 38536 44790 38548
rect 46106 38536 46112 38548
rect 44784 38508 46112 38536
rect 44784 38496 44790 38508
rect 46106 38496 46112 38508
rect 46164 38496 46170 38548
rect 46290 38536 46296 38548
rect 46251 38508 46296 38536
rect 46290 38496 46296 38508
rect 46348 38496 46354 38548
rect 49513 38539 49571 38545
rect 49513 38505 49525 38539
rect 49559 38536 49571 38539
rect 49970 38536 49976 38548
rect 49559 38508 49976 38536
rect 49559 38505 49571 38508
rect 49513 38499 49571 38505
rect 49970 38496 49976 38508
rect 50028 38496 50034 38548
rect 51626 38536 51632 38548
rect 51587 38508 51632 38536
rect 51626 38496 51632 38508
rect 51684 38496 51690 38548
rect 52178 38496 52184 38548
rect 52236 38536 52242 38548
rect 52641 38539 52699 38545
rect 52641 38536 52653 38539
rect 52236 38508 52653 38536
rect 52236 38496 52242 38508
rect 52641 38505 52653 38508
rect 52687 38505 52699 38539
rect 52641 38499 52699 38505
rect 53009 38539 53067 38545
rect 53009 38505 53021 38539
rect 53055 38536 53067 38539
rect 53282 38536 53288 38548
rect 53055 38508 53288 38536
rect 53055 38505 53067 38508
rect 53009 38499 53067 38505
rect 39666 38468 39672 38480
rect 38396 38440 39672 38468
rect 38746 38400 38752 38412
rect 36832 38372 37872 38400
rect 38707 38372 38752 38400
rect 36449 38335 36507 38341
rect 36449 38301 36461 38335
rect 36495 38301 36507 38335
rect 36449 38295 36507 38301
rect 36630 38292 36636 38344
rect 36688 38332 36694 38344
rect 36832 38341 36860 38372
rect 37844 38344 37872 38372
rect 38746 38360 38752 38372
rect 38804 38360 38810 38412
rect 38856 38409 38884 38440
rect 39666 38428 39672 38440
rect 39724 38428 39730 38480
rect 41386 38468 41414 38496
rect 41690 38468 41696 38480
rect 41386 38440 41696 38468
rect 41690 38428 41696 38440
rect 41748 38468 41754 38480
rect 41748 38440 42472 38468
rect 41748 38428 41754 38440
rect 42444 38412 42472 38440
rect 44358 38428 44364 38480
rect 44416 38468 44422 38480
rect 46198 38468 46204 38480
rect 44416 38440 46204 38468
rect 44416 38428 44422 38440
rect 46198 38428 46204 38440
rect 46256 38428 46262 38480
rect 46382 38428 46388 38480
rect 46440 38468 46446 38480
rect 49050 38468 49056 38480
rect 46440 38440 49056 38468
rect 46440 38428 46446 38440
rect 49050 38428 49056 38440
rect 49108 38428 49114 38480
rect 52656 38468 52684 38499
rect 53282 38496 53288 38508
rect 53340 38496 53346 38548
rect 53650 38536 53656 38548
rect 53611 38508 53656 38536
rect 53650 38496 53656 38508
rect 53708 38496 53714 38548
rect 53561 38471 53619 38477
rect 53561 38468 53573 38471
rect 52656 38440 53573 38468
rect 53561 38437 53573 38440
rect 53607 38437 53619 38471
rect 53561 38431 53619 38437
rect 38841 38403 38899 38409
rect 38841 38369 38853 38403
rect 38887 38369 38899 38403
rect 38841 38363 38899 38369
rect 38933 38403 38991 38409
rect 38933 38369 38945 38403
rect 38979 38400 38991 38403
rect 40034 38400 40040 38412
rect 38979 38372 40040 38400
rect 38979 38369 38991 38372
rect 38933 38363 38991 38369
rect 40034 38360 40040 38372
rect 40092 38360 40098 38412
rect 40405 38403 40463 38409
rect 40405 38369 40417 38403
rect 40451 38400 40463 38403
rect 41325 38403 41383 38409
rect 41325 38400 41337 38403
rect 40451 38372 41337 38400
rect 40451 38369 40463 38372
rect 40405 38363 40463 38369
rect 41325 38369 41337 38372
rect 41371 38369 41383 38403
rect 41325 38363 41383 38369
rect 42426 38360 42432 38412
rect 42484 38400 42490 38412
rect 43901 38403 43959 38409
rect 43901 38400 43913 38403
rect 42484 38372 43913 38400
rect 42484 38360 42490 38372
rect 43901 38369 43913 38372
rect 43947 38369 43959 38403
rect 43901 38363 43959 38369
rect 45186 38360 45192 38412
rect 45244 38400 45250 38412
rect 45281 38403 45339 38409
rect 45281 38400 45293 38403
rect 45244 38372 45293 38400
rect 45244 38360 45250 38372
rect 45281 38369 45293 38372
rect 45327 38369 45339 38403
rect 50157 38403 50215 38409
rect 50157 38400 50169 38403
rect 45281 38363 45339 38369
rect 49436 38372 50169 38400
rect 36817 38335 36875 38341
rect 36688 38304 36781 38332
rect 36688 38292 36694 38304
rect 36817 38301 36829 38335
rect 36863 38301 36875 38335
rect 36817 38295 36875 38301
rect 37274 38292 37280 38344
rect 37332 38332 37338 38344
rect 37461 38335 37519 38341
rect 37461 38332 37473 38335
rect 37332 38304 37473 38332
rect 37332 38292 37338 38304
rect 37461 38301 37473 38304
rect 37507 38301 37519 38335
rect 37826 38332 37832 38344
rect 37787 38304 37832 38332
rect 37461 38295 37519 38301
rect 37826 38292 37832 38304
rect 37884 38292 37890 38344
rect 38657 38335 38715 38341
rect 38657 38301 38669 38335
rect 38703 38301 38715 38335
rect 39850 38332 39856 38344
rect 39811 38304 39856 38332
rect 38657 38295 38715 38301
rect 36722 38264 36728 38276
rect 36683 38236 36728 38264
rect 36722 38224 36728 38236
rect 36780 38224 36786 38276
rect 37550 38224 37556 38276
rect 37608 38264 37614 38276
rect 37645 38267 37703 38273
rect 37645 38264 37657 38267
rect 37608 38236 37657 38264
rect 37608 38224 37614 38236
rect 37645 38233 37657 38236
rect 37691 38233 37703 38267
rect 37645 38227 37703 38233
rect 37737 38267 37795 38273
rect 37737 38233 37749 38267
rect 37783 38264 37795 38267
rect 38470 38264 38476 38276
rect 37783 38236 38476 38264
rect 37783 38233 37795 38236
rect 37737 38227 37795 38233
rect 38470 38224 38476 38236
rect 38528 38224 38534 38276
rect 34848 38168 34928 38196
rect 34848 38156 34854 38168
rect 35894 38156 35900 38208
rect 35952 38196 35958 38208
rect 37001 38199 37059 38205
rect 37001 38196 37013 38199
rect 35952 38168 37013 38196
rect 35952 38156 35958 38168
rect 37001 38165 37013 38168
rect 37047 38165 37059 38199
rect 37001 38159 37059 38165
rect 37090 38156 37096 38208
rect 37148 38196 37154 38208
rect 38013 38199 38071 38205
rect 38013 38196 38025 38199
rect 37148 38168 38025 38196
rect 37148 38156 37154 38168
rect 38013 38165 38025 38168
rect 38059 38165 38071 38199
rect 38672 38196 38700 38295
rect 39850 38292 39856 38304
rect 39908 38292 39914 38344
rect 39942 38292 39948 38344
rect 40000 38332 40006 38344
rect 40313 38335 40371 38341
rect 40313 38332 40325 38335
rect 40000 38304 40325 38332
rect 40000 38292 40006 38304
rect 40313 38301 40325 38304
rect 40359 38301 40371 38335
rect 40678 38332 40684 38344
rect 40639 38304 40684 38332
rect 40313 38295 40371 38301
rect 40678 38292 40684 38304
rect 40736 38292 40742 38344
rect 40773 38335 40831 38341
rect 40773 38301 40785 38335
rect 40819 38301 40831 38335
rect 41506 38332 41512 38344
rect 41467 38304 41512 38332
rect 40773 38295 40831 38301
rect 39022 38224 39028 38276
rect 39080 38264 39086 38276
rect 40037 38267 40095 38273
rect 40037 38264 40049 38267
rect 39080 38236 40049 38264
rect 39080 38224 39086 38236
rect 40037 38233 40049 38236
rect 40083 38233 40095 38267
rect 40788 38264 40816 38295
rect 41506 38292 41512 38304
rect 41564 38292 41570 38344
rect 41785 38335 41843 38341
rect 41785 38301 41797 38335
rect 41831 38332 41843 38335
rect 43257 38335 43315 38341
rect 43257 38332 43269 38335
rect 41831 38304 43269 38332
rect 41831 38301 41843 38304
rect 41785 38295 41843 38301
rect 43257 38301 43269 38304
rect 43303 38301 43315 38335
rect 43441 38335 43499 38341
rect 43441 38332 43453 38335
rect 43257 38295 43315 38301
rect 43364 38304 43453 38332
rect 41598 38264 41604 38276
rect 40037 38227 40095 38233
rect 40328 38236 41604 38264
rect 40328 38208 40356 38236
rect 41598 38224 41604 38236
rect 41656 38224 41662 38276
rect 38930 38196 38936 38208
rect 38672 38168 38936 38196
rect 38013 38159 38071 38165
rect 38930 38156 38936 38168
rect 38988 38156 38994 38208
rect 40310 38156 40316 38208
rect 40368 38156 40374 38208
rect 41230 38156 41236 38208
rect 41288 38196 41294 38208
rect 41693 38199 41751 38205
rect 41693 38196 41705 38199
rect 41288 38168 41705 38196
rect 41288 38156 41294 38168
rect 41693 38165 41705 38168
rect 41739 38165 41751 38199
rect 43364 38196 43392 38304
rect 43441 38301 43453 38304
rect 43487 38301 43499 38335
rect 43441 38295 43499 38301
rect 43625 38335 43683 38341
rect 43625 38301 43637 38335
rect 43671 38332 43683 38335
rect 43729 38332 43944 38334
rect 44450 38332 44456 38344
rect 43671 38306 44456 38332
rect 43671 38304 43757 38306
rect 43916 38304 44456 38306
rect 43671 38301 43683 38304
rect 43625 38295 43683 38301
rect 44450 38292 44456 38304
rect 44508 38292 44514 38344
rect 45005 38335 45063 38341
rect 45005 38301 45017 38335
rect 45051 38332 45063 38335
rect 46014 38332 46020 38344
rect 45051 38304 46020 38332
rect 45051 38301 45063 38304
rect 45005 38295 45063 38301
rect 46014 38292 46020 38304
rect 46072 38332 46078 38344
rect 46382 38332 46388 38344
rect 46072 38304 46388 38332
rect 46072 38292 46078 38304
rect 46382 38292 46388 38304
rect 46440 38292 46446 38344
rect 46569 38335 46627 38341
rect 46569 38310 46581 38335
rect 46492 38301 46581 38310
rect 46615 38301 46627 38335
rect 46492 38295 46627 38301
rect 46658 38329 46716 38335
rect 46658 38322 46670 38329
rect 46704 38322 46716 38329
rect 46492 38282 46612 38295
rect 43530 38264 43536 38276
rect 43491 38236 43536 38264
rect 43530 38224 43536 38236
rect 43588 38224 43594 38276
rect 43714 38224 43720 38276
rect 43772 38273 43778 38276
rect 43772 38267 43801 38273
rect 43789 38233 43801 38267
rect 43772 38227 43801 38233
rect 43772 38224 43778 38227
rect 46290 38224 46296 38276
rect 46348 38264 46354 38276
rect 46492 38264 46520 38282
rect 46658 38270 46664 38322
rect 46716 38270 46722 38322
rect 46750 38292 46756 38344
rect 46808 38341 46814 38344
rect 46808 38332 46816 38341
rect 46808 38304 46853 38332
rect 46808 38295 46816 38304
rect 46808 38292 46814 38295
rect 46934 38292 46940 38344
rect 46992 38332 46998 38344
rect 48317 38335 48375 38341
rect 46992 38304 47037 38332
rect 46992 38292 46998 38304
rect 48317 38301 48329 38335
rect 48363 38332 48375 38335
rect 48406 38332 48412 38344
rect 48363 38304 48412 38332
rect 48363 38301 48375 38304
rect 48317 38295 48375 38301
rect 48406 38292 48412 38304
rect 48464 38292 48470 38344
rect 48501 38335 48559 38341
rect 48501 38301 48513 38335
rect 48547 38332 48559 38335
rect 48866 38332 48872 38344
rect 48547 38304 48872 38332
rect 48547 38301 48559 38304
rect 48501 38295 48559 38301
rect 48866 38292 48872 38304
rect 48924 38292 48930 38344
rect 49436 38341 49464 38372
rect 50157 38369 50169 38372
rect 50203 38400 50215 38403
rect 51074 38400 51080 38412
rect 50203 38372 51080 38400
rect 50203 38369 50215 38372
rect 50157 38363 50215 38369
rect 51074 38360 51080 38372
rect 51132 38360 51138 38412
rect 53742 38400 53748 38412
rect 52656 38372 53748 38400
rect 49421 38335 49479 38341
rect 49421 38301 49433 38335
rect 49467 38301 49479 38335
rect 49421 38295 49479 38301
rect 49605 38335 49663 38341
rect 49605 38301 49617 38335
rect 49651 38301 49663 38335
rect 49605 38295 49663 38301
rect 47486 38264 47492 38276
rect 46348 38236 46520 38264
rect 47447 38236 47492 38264
rect 46348 38224 46354 38236
rect 47486 38224 47492 38236
rect 47544 38224 47550 38276
rect 49620 38264 49648 38295
rect 49694 38292 49700 38344
rect 49752 38332 49758 38344
rect 52656 38341 52684 38372
rect 53742 38360 53748 38372
rect 53800 38360 53806 38412
rect 56321 38403 56379 38409
rect 56321 38369 56333 38403
rect 56367 38400 56379 38403
rect 56594 38400 56600 38412
rect 56367 38372 56600 38400
rect 56367 38369 56379 38372
rect 56321 38363 56379 38369
rect 56594 38360 56600 38372
rect 56652 38360 56658 38412
rect 57882 38400 57888 38412
rect 57843 38372 57888 38400
rect 57882 38360 57888 38372
rect 57940 38360 57946 38412
rect 50433 38335 50491 38341
rect 50433 38332 50445 38335
rect 49752 38304 50445 38332
rect 49752 38292 49758 38304
rect 50433 38301 50445 38304
rect 50479 38301 50491 38335
rect 50433 38295 50491 38301
rect 52641 38335 52699 38341
rect 52641 38301 52653 38335
rect 52687 38301 52699 38335
rect 52641 38295 52699 38301
rect 52825 38335 52883 38341
rect 52825 38301 52837 38335
rect 52871 38332 52883 38335
rect 53006 38332 53012 38344
rect 52871 38304 53012 38332
rect 52871 38301 52883 38304
rect 52825 38295 52883 38301
rect 53006 38292 53012 38304
rect 53064 38332 53070 38344
rect 53469 38335 53527 38341
rect 53469 38332 53481 38335
rect 53064 38304 53481 38332
rect 53064 38292 53070 38304
rect 53469 38301 53481 38304
rect 53515 38301 53527 38335
rect 53469 38295 53527 38301
rect 50706 38264 50712 38276
rect 49620 38236 50712 38264
rect 50706 38224 50712 38236
rect 50764 38224 50770 38276
rect 51442 38264 51448 38276
rect 51403 38236 51448 38264
rect 51442 38224 51448 38236
rect 51500 38224 51506 38276
rect 51534 38224 51540 38276
rect 51592 38264 51598 38276
rect 51645 38267 51703 38273
rect 51645 38264 51657 38267
rect 51592 38236 51657 38264
rect 51592 38224 51598 38236
rect 51645 38233 51657 38236
rect 51691 38233 51703 38267
rect 51645 38227 51703 38233
rect 56505 38267 56563 38273
rect 56505 38233 56517 38267
rect 56551 38264 56563 38267
rect 57330 38264 57336 38276
rect 56551 38236 57336 38264
rect 56551 38233 56563 38236
rect 56505 38227 56563 38233
rect 57330 38224 57336 38236
rect 57388 38224 57394 38276
rect 44818 38196 44824 38208
rect 43364 38168 44824 38196
rect 41693 38159 41751 38165
rect 44818 38156 44824 38168
rect 44876 38156 44882 38208
rect 46198 38156 46204 38208
rect 46256 38196 46262 38208
rect 47581 38199 47639 38205
rect 47581 38196 47593 38199
rect 46256 38168 47593 38196
rect 46256 38156 46262 38168
rect 47581 38165 47593 38168
rect 47627 38165 47639 38199
rect 47581 38159 47639 38165
rect 48314 38156 48320 38208
rect 48372 38196 48378 38208
rect 48409 38199 48467 38205
rect 48409 38196 48421 38199
rect 48372 38168 48421 38196
rect 48372 38156 48378 38168
rect 48409 38165 48421 38168
rect 48455 38165 48467 38199
rect 48409 38159 48467 38165
rect 51813 38199 51871 38205
rect 51813 38165 51825 38199
rect 51859 38196 51871 38199
rect 56778 38196 56784 38208
rect 51859 38168 56784 38196
rect 51859 38165 51871 38168
rect 51813 38159 51871 38165
rect 56778 38156 56784 38168
rect 56836 38156 56842 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 22005 37995 22063 38001
rect 22005 37961 22017 37995
rect 22051 37992 22063 37995
rect 22462 37992 22468 38004
rect 22051 37964 22468 37992
rect 22051 37961 22063 37964
rect 22005 37955 22063 37961
rect 22462 37952 22468 37964
rect 22520 37952 22526 38004
rect 22646 37992 22652 38004
rect 22607 37964 22652 37992
rect 22646 37952 22652 37964
rect 22704 37952 22710 38004
rect 23109 37995 23167 38001
rect 23109 37961 23121 37995
rect 23155 37992 23167 37995
rect 24578 37992 24584 38004
rect 23155 37964 24584 37992
rect 23155 37961 23167 37964
rect 23109 37955 23167 37961
rect 24578 37952 24584 37964
rect 24636 37952 24642 38004
rect 24670 37952 24676 38004
rect 24728 37992 24734 38004
rect 24857 37995 24915 38001
rect 24728 37964 24773 37992
rect 24728 37952 24734 37964
rect 24857 37961 24869 37995
rect 24903 37992 24915 37995
rect 25517 37995 25575 38001
rect 25517 37992 25529 37995
rect 24903 37964 25529 37992
rect 24903 37961 24915 37964
rect 24857 37955 24915 37961
rect 25517 37961 25529 37964
rect 25563 37961 25575 37995
rect 26970 37992 26976 38004
rect 25517 37955 25575 37961
rect 25608 37964 26976 37992
rect 25317 37927 25375 37933
rect 21008 37896 23704 37924
rect 20073 37859 20131 37865
rect 20073 37825 20085 37859
rect 20119 37856 20131 37859
rect 20714 37856 20720 37868
rect 20119 37828 20720 37856
rect 20119 37825 20131 37828
rect 20073 37819 20131 37825
rect 20714 37816 20720 37828
rect 20772 37856 20778 37868
rect 21008 37865 21036 37896
rect 20993 37859 21051 37865
rect 20993 37856 21005 37859
rect 20772 37828 21005 37856
rect 20772 37816 20778 37828
rect 20993 37825 21005 37828
rect 21039 37825 21051 37859
rect 22465 37859 22523 37865
rect 22465 37856 22477 37859
rect 20993 37819 21051 37825
rect 22066 37828 22477 37856
rect 20165 37791 20223 37797
rect 20165 37757 20177 37791
rect 20211 37788 20223 37791
rect 20530 37788 20536 37800
rect 20211 37760 20536 37788
rect 20211 37757 20223 37760
rect 20165 37751 20223 37757
rect 20530 37748 20536 37760
rect 20588 37788 20594 37800
rect 22066 37788 22094 37828
rect 22465 37825 22477 37828
rect 22511 37856 22523 37859
rect 23569 37859 23627 37865
rect 23569 37856 23581 37859
rect 22511 37828 23581 37856
rect 22511 37825 22523 37828
rect 22465 37819 22523 37825
rect 23569 37825 23581 37828
rect 23615 37825 23627 37859
rect 23569 37819 23627 37825
rect 22370 37788 22376 37800
rect 20588 37760 22094 37788
rect 22331 37760 22376 37788
rect 20588 37748 20594 37760
rect 22370 37748 22376 37760
rect 22428 37748 22434 37800
rect 22646 37748 22652 37800
rect 22704 37788 22710 37800
rect 22922 37788 22928 37800
rect 22704 37760 22928 37788
rect 22704 37748 22710 37760
rect 22922 37748 22928 37760
rect 22980 37788 22986 37800
rect 23293 37791 23351 37797
rect 23293 37788 23305 37791
rect 22980 37760 23305 37788
rect 22980 37748 22986 37760
rect 23293 37757 23305 37760
rect 23339 37757 23351 37791
rect 23293 37751 23351 37757
rect 23385 37791 23443 37797
rect 23385 37757 23397 37791
rect 23431 37757 23443 37791
rect 23385 37751 23443 37757
rect 23477 37791 23535 37797
rect 23477 37757 23489 37791
rect 23523 37788 23535 37791
rect 23676 37788 23704 37896
rect 25317 37893 25329 37927
rect 25363 37924 25375 37927
rect 25608 37924 25636 37964
rect 26970 37952 26976 37964
rect 27028 37992 27034 38004
rect 28166 37992 28172 38004
rect 27028 37964 28172 37992
rect 27028 37952 27034 37964
rect 28166 37952 28172 37964
rect 28224 37952 28230 38004
rect 29546 37952 29552 38004
rect 29604 37992 29610 38004
rect 29641 37995 29699 38001
rect 29641 37992 29653 37995
rect 29604 37964 29653 37992
rect 29604 37952 29610 37964
rect 29641 37961 29653 37964
rect 29687 37961 29699 37995
rect 29641 37955 29699 37961
rect 30466 37952 30472 38004
rect 30524 37992 30530 38004
rect 31110 37992 31116 38004
rect 30524 37964 31116 37992
rect 30524 37952 30530 37964
rect 31110 37952 31116 37964
rect 31168 37952 31174 38004
rect 32582 37952 32588 38004
rect 32640 37992 32646 38004
rect 32950 37992 32956 38004
rect 32640 37964 32956 37992
rect 32640 37952 32646 37964
rect 32950 37952 32956 37964
rect 33008 37992 33014 38004
rect 33008 37964 35940 37992
rect 33008 37952 33014 37964
rect 25363 37896 25636 37924
rect 25363 37893 25375 37896
rect 25317 37887 25375 37893
rect 30190 37884 30196 37936
rect 30248 37924 30254 37936
rect 35802 37924 35808 37936
rect 30248 37896 32536 37924
rect 30248 37884 30254 37896
rect 24486 37856 24492 37868
rect 24447 37828 24492 37856
rect 24486 37816 24492 37828
rect 24544 37816 24550 37868
rect 24857 37859 24915 37865
rect 24857 37825 24869 37859
rect 24903 37856 24915 37859
rect 25038 37856 25044 37868
rect 24903 37828 25044 37856
rect 24903 37825 24915 37828
rect 24857 37819 24915 37825
rect 25038 37816 25044 37828
rect 25096 37856 25102 37868
rect 26329 37859 26387 37865
rect 26329 37856 26341 37859
rect 25096 37828 25636 37856
rect 25096 37816 25102 37828
rect 23523 37760 23704 37788
rect 23523 37757 23535 37760
rect 23477 37751 23535 37757
rect 22388 37720 22416 37748
rect 23400 37720 23428 37751
rect 22388 37692 23428 37720
rect 20346 37612 20352 37664
rect 20404 37652 20410 37664
rect 20441 37655 20499 37661
rect 20441 37652 20453 37655
rect 20404 37624 20453 37652
rect 20404 37612 20410 37624
rect 20441 37621 20453 37624
rect 20487 37621 20499 37655
rect 20441 37615 20499 37621
rect 20990 37612 20996 37664
rect 21048 37652 21054 37664
rect 21177 37655 21235 37661
rect 21177 37652 21189 37655
rect 21048 37624 21189 37652
rect 21048 37612 21054 37624
rect 21177 37621 21189 37624
rect 21223 37652 21235 37655
rect 22830 37652 22836 37664
rect 21223 37624 22836 37652
rect 21223 37621 21235 37624
rect 21177 37615 21235 37621
rect 22830 37612 22836 37624
rect 22888 37612 22894 37664
rect 25498 37652 25504 37664
rect 25459 37624 25504 37652
rect 25498 37612 25504 37624
rect 25556 37612 25562 37664
rect 25608 37652 25636 37828
rect 25700 37828 26341 37856
rect 25700 37729 25728 37828
rect 26329 37825 26341 37828
rect 26375 37825 26387 37859
rect 26329 37819 26387 37825
rect 29917 37859 29975 37865
rect 29917 37825 29929 37859
rect 29963 37856 29975 37859
rect 30742 37856 30748 37868
rect 29963 37828 30748 37856
rect 29963 37825 29975 37828
rect 29917 37819 29975 37825
rect 30742 37816 30748 37828
rect 30800 37816 30806 37868
rect 32508 37865 32536 37896
rect 34431 37896 35808 37924
rect 32493 37859 32551 37865
rect 32493 37825 32505 37859
rect 32539 37856 32551 37859
rect 33505 37859 33563 37865
rect 33505 37856 33517 37859
rect 32539 37828 33517 37856
rect 32539 37825 32551 37828
rect 32493 37819 32551 37825
rect 33505 37825 33517 37828
rect 33551 37856 33563 37859
rect 34146 37856 34152 37868
rect 33551 37828 34152 37856
rect 33551 37825 33563 37828
rect 33505 37819 33563 37825
rect 34146 37816 34152 37828
rect 34204 37816 34210 37868
rect 29825 37791 29883 37797
rect 29825 37757 29837 37791
rect 29871 37757 29883 37791
rect 30006 37788 30012 37800
rect 29967 37760 30012 37788
rect 29825 37751 29883 37757
rect 25685 37723 25743 37729
rect 25685 37689 25697 37723
rect 25731 37689 25743 37723
rect 26234 37720 26240 37732
rect 25685 37683 25743 37689
rect 25792 37692 26240 37720
rect 25792 37652 25820 37692
rect 26234 37680 26240 37692
rect 26292 37680 26298 37732
rect 29840 37720 29868 37751
rect 30006 37748 30012 37760
rect 30064 37748 30070 37800
rect 30098 37748 30104 37800
rect 30156 37788 30162 37800
rect 31018 37788 31024 37800
rect 30156 37760 30201 37788
rect 30979 37760 31024 37788
rect 30156 37748 30162 37760
rect 31018 37748 31024 37760
rect 31076 37748 31082 37800
rect 32401 37791 32459 37797
rect 32401 37757 32413 37791
rect 32447 37757 32459 37791
rect 32582 37788 32588 37800
rect 32543 37760 32588 37788
rect 32401 37751 32459 37757
rect 31294 37720 31300 37732
rect 29840 37692 31300 37720
rect 31294 37680 31300 37692
rect 31352 37680 31358 37732
rect 32416 37720 32444 37751
rect 32582 37748 32588 37760
rect 32640 37748 32646 37800
rect 32677 37791 32735 37797
rect 32677 37757 32689 37791
rect 32723 37788 32735 37791
rect 33134 37788 33140 37800
rect 32723 37760 33140 37788
rect 32723 37757 32735 37760
rect 32677 37751 32735 37757
rect 33134 37748 33140 37760
rect 33192 37748 33198 37800
rect 33229 37791 33287 37797
rect 33229 37757 33241 37791
rect 33275 37788 33287 37791
rect 33318 37788 33324 37800
rect 33275 37760 33324 37788
rect 33275 37757 33287 37760
rect 33229 37751 33287 37757
rect 33318 37748 33324 37760
rect 33376 37788 33382 37800
rect 34431 37788 34459 37896
rect 35802 37884 35808 37896
rect 35860 37884 35866 37936
rect 34793 37859 34851 37865
rect 34793 37825 34805 37859
rect 34839 37856 34851 37859
rect 35710 37856 35716 37868
rect 34839 37828 35716 37856
rect 34839 37825 34851 37828
rect 34793 37819 34851 37825
rect 35710 37816 35716 37828
rect 35768 37816 35774 37868
rect 33376 37760 34459 37788
rect 34517 37791 34575 37797
rect 33376 37748 33382 37760
rect 34517 37757 34529 37791
rect 34563 37757 34575 37791
rect 34517 37751 34575 37757
rect 33778 37720 33784 37732
rect 32416 37692 33784 37720
rect 33778 37680 33784 37692
rect 33836 37680 33842 37732
rect 26142 37652 26148 37664
rect 25608 37624 25820 37652
rect 26103 37624 26148 37652
rect 26142 37612 26148 37624
rect 26200 37612 26206 37664
rect 32217 37655 32275 37661
rect 32217 37621 32229 37655
rect 32263 37652 32275 37655
rect 34054 37652 34060 37664
rect 32263 37624 34060 37652
rect 32263 37621 32275 37624
rect 32217 37615 32275 37621
rect 34054 37612 34060 37624
rect 34112 37612 34118 37664
rect 34146 37612 34152 37664
rect 34204 37652 34210 37664
rect 34532 37652 34560 37751
rect 35912 37720 35940 37964
rect 36262 37952 36268 38004
rect 36320 37992 36326 38004
rect 39574 37992 39580 38004
rect 36320 37964 39580 37992
rect 36320 37952 36326 37964
rect 39574 37952 39580 37964
rect 39632 37952 39638 38004
rect 39942 37992 39948 38004
rect 39903 37964 39948 37992
rect 39942 37952 39948 37964
rect 40000 37952 40006 38004
rect 41230 37992 41236 38004
rect 41191 37964 41236 37992
rect 41230 37952 41236 37964
rect 41288 37952 41294 38004
rect 42521 37995 42579 38001
rect 42521 37992 42533 37995
rect 41340 37964 42533 37992
rect 36357 37927 36415 37933
rect 36357 37893 36369 37927
rect 36403 37924 36415 37927
rect 36630 37924 36636 37936
rect 36403 37896 36636 37924
rect 36403 37893 36415 37896
rect 36357 37887 36415 37893
rect 36630 37884 36636 37896
rect 36688 37884 36694 37936
rect 37826 37924 37832 37936
rect 37568 37896 37832 37924
rect 36170 37816 36176 37868
rect 36228 37865 36234 37868
rect 36228 37859 36251 37865
rect 36239 37856 36251 37859
rect 36446 37856 36452 37868
rect 36239 37828 36308 37856
rect 36407 37828 36452 37856
rect 36239 37825 36251 37828
rect 36228 37819 36251 37825
rect 36228 37816 36234 37819
rect 36280 37788 36308 37828
rect 36446 37816 36452 37828
rect 36504 37816 36510 37868
rect 37568 37865 37596 37896
rect 37826 37884 37832 37896
rect 37884 37924 37890 37936
rect 37884 37896 38976 37924
rect 37884 37884 37890 37896
rect 38948 37865 38976 37896
rect 39482 37884 39488 37936
rect 39540 37924 39546 37936
rect 39758 37924 39764 37936
rect 39540 37896 39764 37924
rect 39540 37884 39546 37896
rect 39758 37884 39764 37896
rect 39816 37924 39822 37936
rect 40678 37924 40684 37936
rect 39816 37896 40684 37924
rect 39816 37884 39822 37896
rect 40678 37884 40684 37896
rect 40736 37884 40742 37936
rect 41138 37884 41144 37936
rect 41196 37924 41202 37936
rect 41340 37924 41368 37964
rect 42521 37961 42533 37964
rect 42567 37961 42579 37995
rect 42521 37955 42579 37961
rect 43530 37952 43536 38004
rect 43588 37992 43594 38004
rect 43993 37995 44051 38001
rect 43993 37992 44005 37995
rect 43588 37964 44005 37992
rect 43588 37952 43594 37964
rect 43993 37961 44005 37964
rect 44039 37961 44051 37995
rect 43993 37955 44051 37961
rect 45370 37952 45376 38004
rect 45428 37992 45434 38004
rect 45741 37995 45799 38001
rect 45741 37992 45753 37995
rect 45428 37964 45753 37992
rect 45428 37952 45434 37964
rect 45741 37961 45753 37964
rect 45787 37992 45799 37995
rect 46750 37992 46756 38004
rect 45787 37964 46756 37992
rect 45787 37961 45799 37964
rect 45741 37955 45799 37961
rect 46750 37952 46756 37964
rect 46808 37952 46814 38004
rect 47118 37952 47124 38004
rect 47176 37992 47182 38004
rect 48961 37995 49019 38001
rect 48961 37992 48973 37995
rect 47176 37964 48973 37992
rect 47176 37952 47182 37964
rect 47780 37933 47808 37964
rect 48961 37961 48973 37964
rect 49007 37992 49019 37995
rect 49694 37992 49700 38004
rect 49007 37964 49700 37992
rect 49007 37961 49019 37964
rect 48961 37955 49019 37961
rect 49694 37952 49700 37964
rect 49752 37952 49758 38004
rect 52178 37992 52184 38004
rect 52139 37964 52184 37992
rect 52178 37952 52184 37964
rect 52236 37952 52242 38004
rect 43625 37927 43683 37933
rect 41196 37896 41368 37924
rect 41432 37896 43576 37924
rect 41196 37884 41202 37896
rect 36541 37859 36599 37865
rect 36541 37825 36553 37859
rect 36587 37856 36599 37859
rect 37553 37859 37611 37865
rect 37553 37856 37565 37859
rect 36587 37828 37565 37856
rect 36587 37825 36599 37828
rect 36541 37819 36599 37825
rect 37553 37825 37565 37828
rect 37599 37825 37611 37859
rect 37553 37819 37611 37825
rect 38565 37859 38623 37865
rect 38565 37825 38577 37859
rect 38611 37825 38623 37859
rect 38565 37819 38623 37825
rect 38749 37859 38807 37865
rect 38749 37825 38761 37859
rect 38795 37825 38807 37859
rect 38749 37819 38807 37825
rect 38841 37859 38899 37865
rect 38841 37825 38853 37859
rect 38887 37825 38899 37859
rect 38841 37819 38899 37825
rect 38933 37859 38991 37865
rect 38933 37825 38945 37859
rect 38979 37825 38991 37859
rect 40126 37856 40132 37868
rect 40087 37828 40132 37856
rect 38933 37819 38991 37825
rect 37182 37788 37188 37800
rect 36280 37760 37188 37788
rect 37182 37748 37188 37760
rect 37240 37748 37246 37800
rect 37277 37791 37335 37797
rect 37277 37757 37289 37791
rect 37323 37788 37335 37791
rect 37366 37788 37372 37800
rect 37323 37760 37372 37788
rect 37323 37757 37335 37760
rect 37277 37751 37335 37757
rect 37366 37748 37372 37760
rect 37424 37748 37430 37800
rect 38580 37788 38608 37819
rect 37476 37760 38608 37788
rect 37476 37720 37504 37760
rect 35912 37692 37504 37720
rect 37550 37680 37556 37732
rect 37608 37720 37614 37732
rect 38764 37720 38792 37819
rect 37608 37692 38792 37720
rect 38856 37720 38884 37819
rect 40126 37816 40132 37828
rect 40184 37816 40190 37868
rect 40221 37859 40279 37865
rect 40221 37825 40233 37859
rect 40267 37856 40279 37859
rect 40310 37856 40316 37868
rect 40267 37828 40316 37856
rect 40267 37825 40279 37828
rect 40221 37819 40279 37825
rect 40310 37816 40316 37828
rect 40368 37816 40374 37868
rect 40402 37816 40408 37868
rect 40460 37856 40466 37868
rect 41432 37865 41460 37896
rect 43548 37868 43576 37896
rect 43625 37893 43637 37927
rect 43671 37924 43683 37927
rect 44453 37927 44511 37933
rect 44453 37924 44465 37927
rect 43671 37896 44465 37924
rect 43671 37893 43683 37896
rect 43625 37887 43683 37893
rect 44453 37893 44465 37896
rect 44499 37893 44511 37927
rect 44453 37887 44511 37893
rect 47765 37927 47823 37933
rect 47765 37893 47777 37927
rect 47811 37893 47823 37927
rect 47765 37887 47823 37893
rect 50706 37884 50712 37936
rect 50764 37924 50770 37936
rect 51813 37927 51871 37933
rect 51813 37924 51825 37927
rect 50764 37896 51825 37924
rect 50764 37884 50770 37896
rect 51813 37893 51825 37896
rect 51859 37893 51871 37927
rect 51813 37887 51871 37893
rect 51902 37884 51908 37936
rect 51960 37924 51966 37936
rect 52013 37927 52071 37933
rect 52013 37924 52025 37927
rect 51960 37896 52025 37924
rect 51960 37884 51966 37896
rect 52013 37893 52025 37896
rect 52059 37893 52071 37927
rect 52013 37887 52071 37893
rect 40497 37859 40555 37865
rect 40497 37856 40509 37859
rect 40460 37828 40509 37856
rect 40460 37816 40466 37828
rect 40497 37825 40509 37828
rect 40543 37825 40555 37859
rect 40497 37819 40555 37825
rect 41417 37859 41475 37865
rect 41417 37825 41429 37859
rect 41463 37825 41475 37859
rect 41417 37819 41475 37825
rect 41509 37859 41567 37865
rect 41509 37825 41521 37859
rect 41555 37856 41567 37859
rect 41598 37856 41604 37868
rect 41555 37828 41604 37856
rect 41555 37825 41567 37828
rect 41509 37819 41567 37825
rect 41598 37816 41604 37828
rect 41656 37816 41662 37868
rect 41785 37859 41843 37865
rect 41785 37825 41797 37859
rect 41831 37856 41843 37859
rect 42058 37856 42064 37868
rect 41831 37828 42064 37856
rect 41831 37825 41843 37828
rect 41785 37819 41843 37825
rect 42058 37816 42064 37828
rect 42116 37816 42122 37868
rect 42426 37856 42432 37868
rect 42387 37828 42432 37856
rect 42426 37816 42432 37828
rect 42484 37816 42490 37868
rect 42705 37859 42763 37865
rect 42705 37825 42717 37859
rect 42751 37856 42763 37859
rect 42794 37856 42800 37868
rect 42751 37828 42800 37856
rect 42751 37825 42763 37828
rect 42705 37819 42763 37825
rect 42794 37816 42800 37828
rect 42852 37816 42858 37868
rect 43530 37816 43536 37868
rect 43588 37816 43594 37868
rect 43798 37859 43856 37865
rect 43798 37825 43810 37859
rect 43844 37825 43856 37859
rect 43798 37819 43856 37825
rect 44637 37859 44695 37865
rect 44637 37825 44649 37859
rect 44683 37856 44695 37859
rect 45554 37856 45560 37868
rect 44683 37828 45560 37856
rect 44683 37825 44695 37828
rect 44637 37819 44695 37825
rect 41693 37791 41751 37797
rect 41693 37757 41705 37791
rect 41739 37788 41751 37791
rect 42150 37788 42156 37800
rect 41739 37760 42156 37788
rect 41739 37757 41751 37760
rect 41693 37751 41751 37757
rect 42150 37748 42156 37760
rect 42208 37748 42214 37800
rect 43824 37720 43852 37819
rect 45554 37816 45560 37828
rect 45612 37816 45618 37868
rect 46106 37816 46112 37868
rect 46164 37856 46170 37868
rect 46293 37859 46351 37865
rect 46293 37856 46305 37859
rect 46164 37828 46305 37856
rect 46164 37816 46170 37828
rect 46293 37825 46305 37828
rect 46339 37825 46351 37859
rect 46474 37856 46480 37868
rect 46435 37828 46480 37856
rect 46293 37819 46351 37825
rect 46474 37816 46480 37828
rect 46532 37816 46538 37868
rect 47210 37816 47216 37868
rect 47268 37856 47274 37868
rect 47581 37859 47639 37865
rect 47581 37856 47593 37859
rect 47268 37828 47593 37856
rect 47268 37816 47274 37828
rect 47581 37825 47593 37828
rect 47627 37825 47639 37859
rect 47581 37819 47639 37825
rect 47670 37816 47676 37868
rect 47728 37856 47734 37868
rect 48590 37856 48596 37868
rect 47728 37828 48596 37856
rect 47728 37816 47734 37828
rect 48590 37816 48596 37828
rect 48648 37816 48654 37868
rect 48777 37859 48835 37865
rect 48777 37825 48789 37859
rect 48823 37825 48835 37859
rect 48777 37819 48835 37825
rect 48869 37859 48927 37865
rect 48869 37825 48881 37859
rect 48915 37856 48927 37859
rect 49050 37856 49056 37868
rect 48915 37828 49056 37856
rect 48915 37825 48927 37828
rect 48869 37819 48927 37825
rect 44726 37748 44732 37800
rect 44784 37788 44790 37800
rect 44821 37791 44879 37797
rect 44821 37788 44833 37791
rect 44784 37760 44833 37788
rect 44784 37748 44790 37760
rect 44821 37757 44833 37760
rect 44867 37757 44879 37791
rect 44821 37751 44879 37757
rect 44913 37791 44971 37797
rect 44913 37757 44925 37791
rect 44959 37788 44971 37791
rect 45830 37788 45836 37800
rect 44959 37760 45836 37788
rect 44959 37757 44971 37760
rect 44913 37751 44971 37757
rect 45830 37748 45836 37760
rect 45888 37748 45894 37800
rect 46017 37791 46075 37797
rect 46017 37757 46029 37791
rect 46063 37788 46075 37791
rect 46198 37788 46204 37800
rect 46063 37760 46204 37788
rect 46063 37757 46075 37760
rect 46017 37751 46075 37757
rect 46198 37748 46204 37760
rect 46256 37748 46262 37800
rect 46382 37748 46388 37800
rect 46440 37788 46446 37800
rect 48792 37788 48820 37819
rect 49050 37816 49056 37828
rect 49108 37856 49114 37868
rect 49510 37856 49516 37868
rect 49108 37828 49516 37856
rect 49108 37816 49114 37828
rect 49510 37816 49516 37828
rect 49568 37816 49574 37868
rect 49786 37856 49792 37868
rect 49747 37828 49792 37856
rect 49786 37816 49792 37828
rect 49844 37816 49850 37868
rect 49970 37856 49976 37868
rect 49931 37828 49976 37856
rect 49970 37816 49976 37828
rect 50028 37816 50034 37868
rect 50062 37816 50068 37868
rect 50120 37856 50126 37868
rect 50120 37828 50165 37856
rect 50120 37816 50126 37828
rect 50246 37816 50252 37868
rect 50304 37856 50310 37868
rect 50614 37856 50620 37868
rect 50304 37828 50620 37856
rect 50304 37816 50310 37828
rect 50614 37816 50620 37828
rect 50672 37856 50678 37868
rect 50801 37859 50859 37865
rect 50801 37856 50813 37859
rect 50672 37828 50813 37856
rect 50672 37816 50678 37828
rect 50801 37825 50813 37828
rect 50847 37825 50859 37859
rect 50801 37819 50859 37825
rect 52178 37816 52184 37868
rect 52236 37856 52242 37868
rect 53101 37859 53159 37865
rect 53101 37856 53113 37859
rect 52236 37828 53113 37856
rect 52236 37816 52242 37828
rect 53101 37825 53113 37828
rect 53147 37825 53159 37859
rect 56778 37856 56784 37868
rect 56739 37828 56784 37856
rect 53101 37819 53159 37825
rect 56778 37816 56784 37828
rect 56836 37816 56842 37868
rect 46440 37760 48820 37788
rect 46440 37748 46446 37760
rect 49878 37748 49884 37800
rect 49936 37788 49942 37800
rect 50525 37791 50583 37797
rect 50525 37788 50537 37791
rect 49936 37760 50537 37788
rect 49936 37748 49942 37760
rect 50525 37757 50537 37760
rect 50571 37788 50583 37791
rect 53190 37788 53196 37800
rect 50571 37760 51074 37788
rect 53151 37760 53196 37788
rect 50571 37757 50583 37760
rect 50525 37751 50583 37757
rect 45646 37720 45652 37732
rect 38856 37692 45652 37720
rect 37608 37680 37614 37692
rect 45646 37680 45652 37692
rect 45704 37680 45710 37732
rect 46109 37723 46167 37729
rect 46109 37689 46121 37723
rect 46155 37720 46167 37723
rect 47394 37720 47400 37732
rect 46155 37692 47400 37720
rect 46155 37689 46167 37692
rect 46109 37683 46167 37689
rect 47394 37680 47400 37692
rect 47452 37680 47458 37732
rect 48593 37723 48651 37729
rect 48593 37689 48605 37723
rect 48639 37720 48651 37723
rect 48866 37720 48872 37732
rect 48639 37692 48872 37720
rect 48639 37689 48651 37692
rect 48593 37683 48651 37689
rect 48866 37680 48872 37692
rect 48924 37680 48930 37732
rect 49145 37723 49203 37729
rect 49145 37689 49157 37723
rect 49191 37720 49203 37723
rect 50614 37720 50620 37732
rect 49191 37692 50620 37720
rect 49191 37689 49203 37692
rect 49145 37683 49203 37689
rect 50614 37680 50620 37692
rect 50672 37680 50678 37732
rect 36722 37652 36728 37664
rect 34204 37624 34560 37652
rect 36683 37624 36728 37652
rect 34204 37612 34210 37624
rect 36722 37612 36728 37624
rect 36780 37612 36786 37664
rect 37458 37612 37464 37664
rect 37516 37652 37522 37664
rect 39117 37655 39175 37661
rect 39117 37652 39129 37655
rect 37516 37624 39129 37652
rect 37516 37612 37522 37624
rect 39117 37621 39129 37624
rect 39163 37621 39175 37655
rect 39117 37615 39175 37621
rect 40405 37655 40463 37661
rect 40405 37621 40417 37655
rect 40451 37652 40463 37655
rect 41046 37652 41052 37664
rect 40451 37624 41052 37652
rect 40451 37621 40463 37624
rect 40405 37615 40463 37621
rect 41046 37612 41052 37624
rect 41104 37612 41110 37664
rect 46201 37655 46259 37661
rect 46201 37621 46213 37655
rect 46247 37652 46259 37655
rect 47854 37652 47860 37664
rect 46247 37624 47860 37652
rect 46247 37621 46259 37624
rect 46201 37615 46259 37621
rect 47854 37612 47860 37624
rect 47912 37612 47918 37664
rect 47949 37655 48007 37661
rect 47949 37621 47961 37655
rect 47995 37652 48007 37655
rect 48130 37652 48136 37664
rect 47995 37624 48136 37652
rect 47995 37621 48007 37624
rect 47949 37615 48007 37621
rect 48130 37612 48136 37624
rect 48188 37612 48194 37664
rect 49789 37655 49847 37661
rect 49789 37621 49801 37655
rect 49835 37652 49847 37655
rect 50154 37652 50160 37664
rect 49835 37624 50160 37652
rect 49835 37621 49847 37624
rect 49789 37615 49847 37621
rect 50154 37612 50160 37624
rect 50212 37612 50218 37664
rect 51046 37652 51074 37760
rect 53190 37748 53196 37760
rect 53248 37748 53254 37800
rect 56870 37788 56876 37800
rect 56831 37760 56876 37788
rect 56870 37748 56876 37760
rect 56928 37748 56934 37800
rect 57146 37788 57152 37800
rect 57107 37760 57152 37788
rect 57146 37748 57152 37760
rect 57204 37748 57210 37800
rect 53469 37723 53527 37729
rect 53469 37689 53481 37723
rect 53515 37720 53527 37723
rect 53926 37720 53932 37732
rect 53515 37692 53932 37720
rect 53515 37689 53527 37692
rect 53469 37683 53527 37689
rect 53926 37680 53932 37692
rect 53984 37680 53990 37732
rect 51997 37655 52055 37661
rect 51997 37652 52009 37655
rect 51046 37624 52009 37652
rect 51997 37621 52009 37624
rect 52043 37621 52055 37655
rect 51997 37615 52055 37621
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 20625 37451 20683 37457
rect 20625 37417 20637 37451
rect 20671 37448 20683 37451
rect 20898 37448 20904 37460
rect 20671 37420 20904 37448
rect 20671 37417 20683 37420
rect 20625 37411 20683 37417
rect 20898 37408 20904 37420
rect 20956 37408 20962 37460
rect 23382 37448 23388 37460
rect 23343 37420 23388 37448
rect 23382 37408 23388 37420
rect 23440 37408 23446 37460
rect 26510 37408 26516 37460
rect 26568 37448 26574 37460
rect 27246 37448 27252 37460
rect 26568 37420 27252 37448
rect 26568 37408 26574 37420
rect 27246 37408 27252 37420
rect 27304 37448 27310 37460
rect 28261 37451 28319 37457
rect 28261 37448 28273 37451
rect 27304 37420 28273 37448
rect 27304 37408 27310 37420
rect 28261 37417 28273 37420
rect 28307 37417 28319 37451
rect 28261 37411 28319 37417
rect 30285 37451 30343 37457
rect 30285 37417 30297 37451
rect 30331 37448 30343 37451
rect 30374 37448 30380 37460
rect 30331 37420 30380 37448
rect 30331 37417 30343 37420
rect 30285 37411 30343 37417
rect 30374 37408 30380 37420
rect 30432 37408 30438 37460
rect 31110 37408 31116 37460
rect 31168 37448 31174 37460
rect 34146 37448 34152 37460
rect 31168 37420 34152 37448
rect 31168 37408 31174 37420
rect 20441 37315 20499 37321
rect 20441 37281 20453 37315
rect 20487 37312 20499 37315
rect 20806 37312 20812 37324
rect 20487 37284 20812 37312
rect 20487 37281 20499 37284
rect 20441 37275 20499 37281
rect 20806 37272 20812 37284
rect 20864 37272 20870 37324
rect 31294 37272 31300 37324
rect 31352 37312 31358 37324
rect 31665 37315 31723 37321
rect 31352 37284 31524 37312
rect 31352 37272 31358 37284
rect 31496 37256 31524 37284
rect 31665 37281 31677 37315
rect 31711 37312 31723 37315
rect 32306 37312 32312 37324
rect 31711 37284 32312 37312
rect 31711 37281 31723 37284
rect 31665 37275 31723 37281
rect 32306 37272 32312 37284
rect 32364 37272 32370 37324
rect 33336 37321 33364 37420
rect 34146 37408 34152 37420
rect 34204 37408 34210 37460
rect 34330 37408 34336 37460
rect 34388 37448 34394 37460
rect 34388 37420 36400 37448
rect 34388 37408 34394 37420
rect 33778 37340 33784 37392
rect 33836 37380 33842 37392
rect 33836 37352 34376 37380
rect 33836 37340 33842 37352
rect 33321 37315 33379 37321
rect 33321 37281 33333 37315
rect 33367 37281 33379 37315
rect 33321 37275 33379 37281
rect 33410 37272 33416 37324
rect 33468 37312 33474 37324
rect 34348 37312 34376 37352
rect 36372 37324 36400 37420
rect 36446 37408 36452 37460
rect 36504 37448 36510 37460
rect 39298 37448 39304 37460
rect 36504 37420 39304 37448
rect 36504 37408 36510 37420
rect 39298 37408 39304 37420
rect 39356 37448 39362 37460
rect 39356 37420 40540 37448
rect 39356 37408 39362 37420
rect 37366 37340 37372 37392
rect 37424 37380 37430 37392
rect 37424 37352 37964 37380
rect 37424 37340 37430 37352
rect 34790 37312 34796 37324
rect 33468 37284 33732 37312
rect 34348 37284 34796 37312
rect 33468 37272 33474 37284
rect 20346 37244 20352 37256
rect 20307 37216 20352 37244
rect 20346 37204 20352 37216
rect 20404 37204 20410 37256
rect 20622 37204 20628 37256
rect 20680 37244 20686 37256
rect 21361 37247 21419 37253
rect 21361 37244 21373 37247
rect 20680 37216 21373 37244
rect 20680 37204 20686 37216
rect 21361 37213 21373 37216
rect 21407 37244 21419 37247
rect 21407 37216 22094 37244
rect 21407 37213 21419 37216
rect 21361 37207 21419 37213
rect 21634 37185 21640 37188
rect 21628 37176 21640 37185
rect 21595 37148 21640 37176
rect 21628 37139 21640 37148
rect 21634 37136 21640 37139
rect 21692 37136 21698 37188
rect 22066 37176 22094 37216
rect 22370 37204 22376 37256
rect 22428 37244 22434 37256
rect 23201 37247 23259 37253
rect 23201 37244 23213 37247
rect 22428 37216 23213 37244
rect 22428 37204 22434 37216
rect 23201 37213 23213 37216
rect 23247 37213 23259 37247
rect 23201 37207 23259 37213
rect 25869 37247 25927 37253
rect 25869 37213 25881 37247
rect 25915 37244 25927 37247
rect 26694 37244 26700 37256
rect 25915 37216 26700 37244
rect 25915 37213 25927 37216
rect 25869 37207 25927 37213
rect 25884 37176 25912 37207
rect 26694 37204 26700 37216
rect 26752 37204 26758 37256
rect 28169 37247 28227 37253
rect 28169 37213 28181 37247
rect 28215 37244 28227 37247
rect 29638 37244 29644 37256
rect 28215 37216 29644 37244
rect 28215 37213 28227 37216
rect 28169 37207 28227 37213
rect 29638 37204 29644 37216
rect 29696 37204 29702 37256
rect 30006 37204 30012 37256
rect 30064 37244 30070 37256
rect 30469 37247 30527 37253
rect 30469 37244 30481 37247
rect 30064 37216 30481 37244
rect 30064 37204 30070 37216
rect 30469 37213 30481 37216
rect 30515 37213 30527 37247
rect 30469 37207 30527 37213
rect 30561 37247 30619 37253
rect 30561 37213 30573 37247
rect 30607 37244 30619 37247
rect 31018 37244 31024 37256
rect 30607 37216 31024 37244
rect 30607 37213 30619 37216
rect 30561 37207 30619 37213
rect 31018 37204 31024 37216
rect 31076 37204 31082 37256
rect 31202 37204 31208 37256
rect 31260 37244 31266 37256
rect 31389 37247 31447 37253
rect 31389 37244 31401 37247
rect 31260 37216 31401 37244
rect 31260 37204 31266 37216
rect 31389 37213 31401 37216
rect 31435 37213 31447 37247
rect 31389 37207 31447 37213
rect 31478 37204 31484 37256
rect 31536 37244 31542 37256
rect 31846 37253 31852 37256
rect 31573 37247 31631 37253
rect 31573 37244 31585 37247
rect 31536 37216 31585 37244
rect 31536 37204 31542 37216
rect 31573 37213 31585 37216
rect 31619 37213 31631 37247
rect 31573 37207 31631 37213
rect 31803 37247 31852 37253
rect 31803 37213 31815 37247
rect 31849 37213 31852 37247
rect 31803 37207 31852 37213
rect 31846 37204 31852 37207
rect 31904 37204 31910 37256
rect 31941 37247 31999 37253
rect 31941 37213 31953 37247
rect 31987 37213 31999 37247
rect 31941 37207 31999 37213
rect 33597 37247 33655 37253
rect 33597 37213 33609 37247
rect 33643 37213 33655 37247
rect 33704 37244 33732 37284
rect 34790 37272 34796 37284
rect 34848 37312 34854 37324
rect 34977 37315 35035 37321
rect 34977 37312 34989 37315
rect 34848 37284 34989 37312
rect 34848 37272 34854 37284
rect 34977 37281 34989 37284
rect 35023 37281 35035 37315
rect 36354 37312 36360 37324
rect 36267 37284 36360 37312
rect 34977 37275 35035 37281
rect 36354 37272 36360 37284
rect 36412 37312 36418 37324
rect 36541 37315 36599 37321
rect 36541 37312 36553 37315
rect 36412 37284 36553 37312
rect 36412 37272 36418 37284
rect 36541 37281 36553 37284
rect 36587 37281 36599 37315
rect 36541 37275 36599 37281
rect 36817 37315 36875 37321
rect 36817 37281 36829 37315
rect 36863 37312 36875 37315
rect 37550 37312 37556 37324
rect 36863 37284 37556 37312
rect 36863 37281 36875 37284
rect 36817 37275 36875 37281
rect 34701 37247 34759 37253
rect 34701 37244 34713 37247
rect 33704 37216 34713 37244
rect 33597 37207 33655 37213
rect 34701 37213 34713 37216
rect 34747 37244 34759 37247
rect 35710 37244 35716 37256
rect 34747 37216 35716 37244
rect 34747 37213 34759 37216
rect 34701 37207 34759 37213
rect 26142 37185 26148 37188
rect 26136 37176 26148 37185
rect 22066 37148 25912 37176
rect 26103 37148 26148 37176
rect 26136 37139 26148 37148
rect 26142 37136 26148 37139
rect 26200 37136 26206 37188
rect 30282 37176 30288 37188
rect 30243 37148 30288 37176
rect 30282 37136 30288 37148
rect 30340 37136 30346 37188
rect 31662 37136 31668 37188
rect 31720 37176 31726 37188
rect 31956 37176 31984 37207
rect 33612 37176 33640 37207
rect 35710 37204 35716 37216
rect 35768 37244 35774 37256
rect 36078 37244 36084 37256
rect 35768 37216 36084 37244
rect 35768 37204 35774 37216
rect 36078 37204 36084 37216
rect 36136 37204 36142 37256
rect 33962 37176 33968 37188
rect 31720 37148 33456 37176
rect 33612 37148 33968 37176
rect 31720 37136 31726 37148
rect 22370 37068 22376 37120
rect 22428 37108 22434 37120
rect 22741 37111 22799 37117
rect 22741 37108 22753 37111
rect 22428 37080 22753 37108
rect 22428 37068 22434 37080
rect 22741 37077 22753 37080
rect 22787 37077 22799 37111
rect 22741 37071 22799 37077
rect 26234 37068 26240 37120
rect 26292 37108 26298 37120
rect 27249 37111 27307 37117
rect 27249 37108 27261 37111
rect 26292 37080 27261 37108
rect 26292 37068 26298 37080
rect 27249 37077 27261 37080
rect 27295 37108 27307 37111
rect 31846 37108 31852 37120
rect 27295 37080 31852 37108
rect 27295 37077 27307 37080
rect 27249 37071 27307 37077
rect 31846 37068 31852 37080
rect 31904 37068 31910 37120
rect 32122 37108 32128 37120
rect 32083 37080 32128 37108
rect 32122 37068 32128 37080
rect 32180 37068 32186 37120
rect 33428 37108 33456 37148
rect 33962 37136 33968 37148
rect 34020 37136 34026 37188
rect 36556 37176 36584 37275
rect 37550 37272 37556 37284
rect 37608 37272 37614 37324
rect 37274 37204 37280 37256
rect 37332 37244 37338 37256
rect 37829 37247 37887 37253
rect 37829 37244 37841 37247
rect 37332 37216 37841 37244
rect 37332 37204 37338 37216
rect 37829 37213 37841 37216
rect 37875 37213 37887 37247
rect 37936 37244 37964 37352
rect 38746 37340 38752 37392
rect 38804 37380 38810 37392
rect 40129 37383 40187 37389
rect 40129 37380 40141 37383
rect 38804 37352 40141 37380
rect 38804 37340 38810 37352
rect 40129 37349 40141 37352
rect 40175 37349 40187 37383
rect 40512 37380 40540 37420
rect 40586 37408 40592 37460
rect 40644 37448 40650 37460
rect 42058 37448 42064 37460
rect 40644 37420 42064 37448
rect 40644 37408 40650 37420
rect 42058 37408 42064 37420
rect 42116 37408 42122 37460
rect 42150 37408 42156 37460
rect 42208 37448 42214 37460
rect 42981 37451 43039 37457
rect 42981 37448 42993 37451
rect 42208 37420 42993 37448
rect 42208 37408 42214 37420
rect 42981 37417 42993 37420
rect 43027 37417 43039 37451
rect 42981 37411 43039 37417
rect 44726 37408 44732 37460
rect 44784 37448 44790 37460
rect 45186 37448 45192 37460
rect 44784 37420 45192 37448
rect 44784 37408 44790 37420
rect 45186 37408 45192 37420
rect 45244 37448 45250 37460
rect 45373 37451 45431 37457
rect 45373 37448 45385 37451
rect 45244 37420 45385 37448
rect 45244 37408 45250 37420
rect 45373 37417 45385 37420
rect 45419 37417 45431 37451
rect 45373 37411 45431 37417
rect 45925 37451 45983 37457
rect 45925 37417 45937 37451
rect 45971 37448 45983 37451
rect 46014 37448 46020 37460
rect 45971 37420 46020 37448
rect 45971 37417 45983 37420
rect 45925 37411 45983 37417
rect 46014 37408 46020 37420
rect 46072 37408 46078 37460
rect 47213 37451 47271 37457
rect 47213 37417 47225 37451
rect 47259 37417 47271 37451
rect 47394 37448 47400 37460
rect 47355 37420 47400 37448
rect 47213 37411 47271 37417
rect 41414 37380 41420 37392
rect 40512 37352 41420 37380
rect 40129 37343 40187 37349
rect 41414 37340 41420 37352
rect 41472 37340 41478 37392
rect 42702 37340 42708 37392
rect 42760 37380 42766 37392
rect 46382 37380 46388 37392
rect 42760 37352 46388 37380
rect 42760 37340 42766 37352
rect 46382 37340 46388 37352
rect 46440 37340 46446 37392
rect 47228 37380 47256 37411
rect 47394 37408 47400 37420
rect 47452 37408 47458 37460
rect 47854 37448 47860 37460
rect 47815 37420 47860 37448
rect 47854 37408 47860 37420
rect 47912 37408 47918 37460
rect 48130 37380 48136 37392
rect 47228 37352 48136 37380
rect 48130 37340 48136 37352
rect 48188 37340 48194 37392
rect 56042 37340 56048 37392
rect 56100 37380 56106 37392
rect 57793 37383 57851 37389
rect 56100 37352 57284 37380
rect 56100 37340 56106 37352
rect 43625 37315 43683 37321
rect 40420 37284 40908 37312
rect 40420 37256 40448 37284
rect 38197 37247 38255 37253
rect 38197 37244 38209 37247
rect 37936 37216 38209 37244
rect 37829 37207 37887 37213
rect 38197 37213 38209 37216
rect 38243 37213 38255 37247
rect 40402 37244 40408 37256
rect 38197 37207 38255 37213
rect 39408 37216 40408 37244
rect 38013 37179 38071 37185
rect 38013 37176 38025 37179
rect 36556 37148 38025 37176
rect 38013 37145 38025 37148
rect 38059 37145 38071 37179
rect 38013 37139 38071 37145
rect 38105 37179 38163 37185
rect 38105 37145 38117 37179
rect 38151 37176 38163 37179
rect 39408 37176 39436 37216
rect 40402 37204 40408 37216
rect 40460 37204 40466 37256
rect 40586 37204 40592 37256
rect 40644 37244 40650 37256
rect 40644 37216 40689 37244
rect 40644 37204 40650 37216
rect 40880 37185 40908 37284
rect 43625 37281 43637 37315
rect 43671 37312 43683 37315
rect 44726 37312 44732 37324
rect 43671 37284 44732 37312
rect 43671 37281 43683 37284
rect 43625 37275 43683 37281
rect 44726 37272 44732 37284
rect 44784 37272 44790 37324
rect 45370 37312 45376 37324
rect 45204 37284 45376 37312
rect 40957 37247 41015 37253
rect 40957 37213 40969 37247
rect 41003 37244 41015 37247
rect 41046 37244 41052 37256
rect 41003 37216 41052 37244
rect 41003 37213 41015 37216
rect 40957 37207 41015 37213
rect 41046 37204 41052 37216
rect 41104 37204 41110 37256
rect 41138 37204 41144 37256
rect 41196 37244 41202 37256
rect 42426 37244 42432 37256
rect 41196 37216 42432 37244
rect 41196 37204 41202 37216
rect 42426 37204 42432 37216
rect 42484 37204 42490 37256
rect 45204 37253 45232 37284
rect 45370 37272 45376 37284
rect 45428 37272 45434 37324
rect 45465 37315 45523 37321
rect 45465 37281 45477 37315
rect 45511 37312 45523 37315
rect 46290 37312 46296 37324
rect 45511 37284 46296 37312
rect 45511 37281 45523 37284
rect 45465 37275 45523 37281
rect 46290 37272 46296 37284
rect 46348 37312 46354 37324
rect 47210 37312 47216 37324
rect 46348 37284 47216 37312
rect 46348 37272 46354 37284
rect 47210 37272 47216 37284
rect 47268 37272 47274 37324
rect 49050 37312 49056 37324
rect 47504 37284 49056 37312
rect 47504 37256 47532 37284
rect 49050 37272 49056 37284
rect 49108 37272 49114 37324
rect 49510 37312 49516 37324
rect 49160 37284 49516 37312
rect 45189 37247 45247 37253
rect 45189 37213 45201 37247
rect 45235 37213 45247 37247
rect 45189 37207 45247 37213
rect 45278 37204 45284 37256
rect 45336 37244 45342 37256
rect 45925 37247 45983 37253
rect 45925 37244 45937 37247
rect 45336 37216 45937 37244
rect 45336 37204 45342 37216
rect 45925 37213 45937 37216
rect 45971 37213 45983 37247
rect 46106 37244 46112 37256
rect 46067 37216 46112 37244
rect 45925 37207 45983 37213
rect 38151 37148 39436 37176
rect 39945 37179 40003 37185
rect 38151 37145 38163 37148
rect 38105 37139 38163 37145
rect 39945 37145 39957 37179
rect 39991 37145 40003 37179
rect 39945 37139 40003 37145
rect 40773 37179 40831 37185
rect 40773 37145 40785 37179
rect 40819 37145 40831 37179
rect 40773 37139 40831 37145
rect 40865 37179 40923 37185
rect 40865 37145 40877 37179
rect 40911 37145 40923 37179
rect 42150 37176 42156 37188
rect 40865 37139 40923 37145
rect 40972 37148 42156 37176
rect 34790 37108 34796 37120
rect 33428 37080 34796 37108
rect 34790 37068 34796 37080
rect 34848 37108 34854 37120
rect 36170 37108 36176 37120
rect 34848 37080 36176 37108
rect 34848 37068 34854 37080
rect 36170 37068 36176 37080
rect 36228 37068 36234 37120
rect 38378 37108 38384 37120
rect 38339 37080 38384 37108
rect 38378 37068 38384 37080
rect 38436 37068 38442 37120
rect 39960 37108 39988 37139
rect 40586 37108 40592 37120
rect 39960 37080 40592 37108
rect 40586 37068 40592 37080
rect 40644 37068 40650 37120
rect 40788 37108 40816 37139
rect 40972 37108 41000 37148
rect 42150 37136 42156 37148
rect 42208 37136 42214 37188
rect 43349 37179 43407 37185
rect 43349 37145 43361 37179
rect 43395 37176 43407 37179
rect 45940 37176 45968 37207
rect 46106 37204 46112 37216
rect 46164 37204 46170 37256
rect 46198 37204 46204 37256
rect 46256 37244 46262 37256
rect 46474 37244 46480 37256
rect 46256 37216 46480 37244
rect 46256 37204 46262 37216
rect 46474 37204 46480 37216
rect 46532 37204 46538 37256
rect 47486 37244 47492 37256
rect 46952 37216 47492 37244
rect 46952 37176 46980 37216
rect 47486 37204 47492 37216
rect 47544 37204 47550 37256
rect 48130 37244 48136 37256
rect 48091 37216 48136 37244
rect 48130 37204 48136 37216
rect 48188 37204 48194 37256
rect 48498 37204 48504 37256
rect 48556 37244 48562 37256
rect 49160 37253 49188 37284
rect 49510 37272 49516 37284
rect 49568 37272 49574 37324
rect 49694 37272 49700 37324
rect 49752 37312 49758 37324
rect 50341 37315 50399 37321
rect 50341 37312 50353 37315
rect 49752 37284 50353 37312
rect 49752 37272 49758 37284
rect 50341 37281 50353 37284
rect 50387 37281 50399 37315
rect 50341 37275 50399 37281
rect 50525 37315 50583 37321
rect 50525 37281 50537 37315
rect 50571 37312 50583 37315
rect 51258 37312 51264 37324
rect 50571 37284 51264 37312
rect 50571 37281 50583 37284
rect 50525 37275 50583 37281
rect 51258 37272 51264 37284
rect 51316 37312 51322 37324
rect 51810 37312 51816 37324
rect 51316 37284 51816 37312
rect 51316 37272 51322 37284
rect 51810 37272 51816 37284
rect 51868 37272 51874 37324
rect 56594 37312 56600 37324
rect 56555 37284 56600 37312
rect 56594 37272 56600 37284
rect 56652 37272 56658 37324
rect 57256 37321 57284 37352
rect 57793 37349 57805 37383
rect 57839 37349 57851 37383
rect 57793 37343 57851 37349
rect 57241 37315 57299 37321
rect 57241 37281 57253 37315
rect 57287 37281 57299 37315
rect 57241 37275 57299 37281
rect 48869 37247 48927 37253
rect 48869 37244 48881 37247
rect 48556 37216 48881 37244
rect 48556 37204 48562 37216
rect 48869 37213 48881 37216
rect 48915 37213 48927 37247
rect 48869 37207 48927 37213
rect 49145 37247 49203 37253
rect 49145 37213 49157 37247
rect 49191 37213 49203 37247
rect 49145 37207 49203 37213
rect 49237 37247 49295 37253
rect 49237 37213 49249 37247
rect 49283 37244 49295 37247
rect 50246 37244 50252 37256
rect 49283 37216 50252 37244
rect 49283 37213 49295 37216
rect 49237 37207 49295 37213
rect 50246 37204 50252 37216
rect 50304 37204 50310 37256
rect 50433 37247 50491 37253
rect 50433 37213 50445 37247
rect 50479 37213 50491 37247
rect 50433 37207 50491 37213
rect 43395 37148 45140 37176
rect 45940 37148 46980 37176
rect 47029 37179 47087 37185
rect 43395 37145 43407 37148
rect 43349 37139 43407 37145
rect 40788 37080 41000 37108
rect 41141 37111 41199 37117
rect 41141 37077 41153 37111
rect 41187 37108 41199 37111
rect 41506 37108 41512 37120
rect 41187 37080 41512 37108
rect 41187 37077 41199 37080
rect 41141 37071 41199 37077
rect 41506 37068 41512 37080
rect 41564 37068 41570 37120
rect 43438 37068 43444 37120
rect 43496 37108 43502 37120
rect 43496 37080 43541 37108
rect 43496 37068 43502 37080
rect 44450 37068 44456 37120
rect 44508 37108 44514 37120
rect 45005 37111 45063 37117
rect 45005 37108 45017 37111
rect 44508 37080 45017 37108
rect 44508 37068 44514 37080
rect 45005 37077 45017 37080
rect 45051 37077 45063 37111
rect 45112 37108 45140 37148
rect 47029 37145 47041 37179
rect 47075 37145 47087 37179
rect 47029 37139 47087 37145
rect 47245 37179 47303 37185
rect 47245 37145 47257 37179
rect 47291 37176 47303 37179
rect 47857 37179 47915 37185
rect 47857 37176 47869 37179
rect 47291 37148 47869 37176
rect 47291 37145 47303 37148
rect 47245 37139 47303 37145
rect 47857 37145 47869 37148
rect 47903 37176 47915 37179
rect 48314 37176 48320 37188
rect 47903 37148 48320 37176
rect 47903 37145 47915 37148
rect 47857 37139 47915 37145
rect 45646 37108 45652 37120
rect 45112 37080 45652 37108
rect 45005 37071 45063 37077
rect 45646 37068 45652 37080
rect 45704 37068 45710 37120
rect 47044 37108 47072 37139
rect 48314 37136 48320 37148
rect 48372 37136 48378 37188
rect 48406 37136 48412 37188
rect 48464 37176 48470 37188
rect 49053 37179 49111 37185
rect 49053 37176 49065 37179
rect 48464 37148 49065 37176
rect 48464 37136 48470 37148
rect 49053 37145 49065 37148
rect 49099 37145 49111 37179
rect 50448 37176 50476 37207
rect 50614 37204 50620 37256
rect 50672 37244 50678 37256
rect 56689 37247 56747 37253
rect 50672 37216 50717 37244
rect 50672 37204 50678 37216
rect 56689 37213 56701 37247
rect 56735 37244 56747 37247
rect 57808 37244 57836 37343
rect 56735 37216 57836 37244
rect 56735 37213 56747 37216
rect 56689 37207 56747 37213
rect 57974 37204 57980 37256
rect 58032 37244 58038 37256
rect 58069 37247 58127 37253
rect 58069 37244 58081 37247
rect 58032 37216 58081 37244
rect 58032 37204 58038 37216
rect 58069 37213 58081 37216
rect 58115 37213 58127 37247
rect 58069 37207 58127 37213
rect 49053 37139 49111 37145
rect 49160 37148 50476 37176
rect 47670 37108 47676 37120
rect 47044 37080 47676 37108
rect 47670 37068 47676 37080
rect 47728 37108 47734 37120
rect 48041 37111 48099 37117
rect 48041 37108 48053 37111
rect 47728 37080 48053 37108
rect 47728 37068 47734 37080
rect 48041 37077 48053 37080
rect 48087 37077 48099 37111
rect 48041 37071 48099 37077
rect 48130 37068 48136 37120
rect 48188 37108 48194 37120
rect 49160 37108 49188 37148
rect 57146 37136 57152 37188
rect 57204 37176 57210 37188
rect 57793 37179 57851 37185
rect 57793 37176 57805 37179
rect 57204 37148 57805 37176
rect 57204 37136 57210 37148
rect 57793 37145 57805 37148
rect 57839 37145 57851 37179
rect 57793 37139 57851 37145
rect 48188 37080 49188 37108
rect 49421 37111 49479 37117
rect 48188 37068 48194 37080
rect 49421 37077 49433 37111
rect 49467 37108 49479 37111
rect 49970 37108 49976 37120
rect 49467 37080 49976 37108
rect 49467 37077 49479 37080
rect 49421 37071 49479 37077
rect 49970 37068 49976 37080
rect 50028 37068 50034 37120
rect 50157 37111 50215 37117
rect 50157 37077 50169 37111
rect 50203 37108 50215 37111
rect 52178 37108 52184 37120
rect 50203 37080 52184 37108
rect 50203 37077 50215 37080
rect 50157 37071 50215 37077
rect 52178 37068 52184 37080
rect 52236 37068 52242 37120
rect 56778 37068 56784 37120
rect 56836 37108 56842 37120
rect 57977 37111 58035 37117
rect 57977 37108 57989 37111
rect 56836 37080 57989 37108
rect 56836 37068 56842 37080
rect 57977 37077 57989 37080
rect 58023 37077 58035 37111
rect 57977 37071 58035 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 23109 36907 23167 36913
rect 23109 36873 23121 36907
rect 23155 36904 23167 36907
rect 24486 36904 24492 36916
rect 23155 36876 24492 36904
rect 23155 36873 23167 36876
rect 23109 36867 23167 36873
rect 24486 36864 24492 36876
rect 24544 36864 24550 36916
rect 31662 36904 31668 36916
rect 24596 36876 31668 36904
rect 22554 36796 22560 36848
rect 22612 36836 22618 36848
rect 24596 36836 24624 36876
rect 31662 36864 31668 36876
rect 31720 36864 31726 36916
rect 31846 36864 31852 36916
rect 31904 36904 31910 36916
rect 32214 36904 32220 36916
rect 31904 36876 32220 36904
rect 31904 36864 31910 36876
rect 32214 36864 32220 36876
rect 32272 36904 32278 36916
rect 32950 36904 32956 36916
rect 32272 36876 32956 36904
rect 32272 36864 32278 36876
rect 32950 36864 32956 36876
rect 33008 36864 33014 36916
rect 33134 36864 33140 36916
rect 33192 36904 33198 36916
rect 33505 36907 33563 36913
rect 33505 36904 33517 36907
rect 33192 36876 33517 36904
rect 33192 36864 33198 36876
rect 33505 36873 33517 36876
rect 33551 36873 33563 36907
rect 44818 36904 44824 36916
rect 33505 36867 33563 36873
rect 33612 36876 44680 36904
rect 44779 36876 44824 36904
rect 22612 36808 24624 36836
rect 28490 36808 29500 36836
rect 22612 36796 22618 36808
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36768 22063 36771
rect 22370 36768 22376 36780
rect 22051 36740 22376 36768
rect 22051 36737 22063 36740
rect 22005 36731 22063 36737
rect 22370 36728 22376 36740
rect 22428 36728 22434 36780
rect 22830 36768 22836 36780
rect 22791 36740 22836 36768
rect 22830 36728 22836 36740
rect 22888 36728 22894 36780
rect 22922 36728 22928 36780
rect 22980 36768 22986 36780
rect 28490 36777 28518 36808
rect 25961 36771 26019 36777
rect 22980 36740 23025 36768
rect 22980 36728 22986 36740
rect 25961 36737 25973 36771
rect 26007 36768 26019 36771
rect 28445 36771 28518 36777
rect 26007 36740 27476 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 22097 36703 22155 36709
rect 22097 36669 22109 36703
rect 22143 36700 22155 36703
rect 22186 36700 22192 36712
rect 22143 36672 22192 36700
rect 22143 36669 22155 36672
rect 22097 36663 22155 36669
rect 22186 36660 22192 36672
rect 22244 36700 22250 36712
rect 23109 36703 23167 36709
rect 23109 36700 23121 36703
rect 22244 36672 23121 36700
rect 22244 36660 22250 36672
rect 23109 36669 23121 36672
rect 23155 36669 23167 36703
rect 23109 36663 23167 36669
rect 26237 36703 26295 36709
rect 26237 36669 26249 36703
rect 26283 36700 26295 36703
rect 26326 36700 26332 36712
rect 26283 36672 26332 36700
rect 26283 36669 26295 36672
rect 26237 36663 26295 36669
rect 26326 36660 26332 36672
rect 26384 36660 26390 36712
rect 27448 36700 27476 36740
rect 28445 36737 28457 36771
rect 28491 36737 28518 36771
rect 29362 36768 29368 36780
rect 29323 36740 29368 36768
rect 28445 36731 28518 36737
rect 28460 36730 28518 36731
rect 29362 36728 29368 36740
rect 29420 36728 29426 36780
rect 29472 36768 29500 36808
rect 29638 36796 29644 36848
rect 29696 36836 29702 36848
rect 31113 36839 31171 36845
rect 31113 36836 31125 36839
rect 29696 36808 31125 36836
rect 29696 36796 29702 36808
rect 31113 36805 31125 36808
rect 31159 36805 31171 36839
rect 31113 36799 31171 36805
rect 32398 36768 32404 36780
rect 29472 36740 32404 36768
rect 32398 36728 32404 36740
rect 32456 36728 32462 36780
rect 33410 36768 33416 36780
rect 33371 36740 33416 36768
rect 33410 36728 33416 36740
rect 33468 36728 33474 36780
rect 33612 36777 33640 36876
rect 34146 36796 34152 36848
rect 34204 36836 34210 36848
rect 35802 36836 35808 36848
rect 34204 36808 34560 36836
rect 34204 36796 34210 36808
rect 33597 36771 33655 36777
rect 33597 36737 33609 36771
rect 33643 36737 33655 36771
rect 33597 36731 33655 36737
rect 33778 36728 33784 36780
rect 33836 36768 33842 36780
rect 34532 36777 34560 36808
rect 35176 36808 35808 36836
rect 34241 36771 34299 36777
rect 34241 36768 34253 36771
rect 33836 36740 34253 36768
rect 33836 36728 33842 36740
rect 34241 36737 34253 36740
rect 34287 36737 34299 36771
rect 34241 36731 34299 36737
rect 34517 36771 34575 36777
rect 34517 36737 34529 36771
rect 34563 36737 34575 36771
rect 34517 36731 34575 36737
rect 27448 36672 28488 36700
rect 22373 36635 22431 36641
rect 22373 36601 22385 36635
rect 22419 36632 22431 36635
rect 23198 36632 23204 36644
rect 22419 36604 23204 36632
rect 22419 36601 22431 36604
rect 22373 36595 22431 36601
rect 23198 36592 23204 36604
rect 23256 36592 23262 36644
rect 28460 36632 28488 36672
rect 28626 36660 28632 36712
rect 28684 36700 28690 36712
rect 28721 36703 28779 36709
rect 28721 36700 28733 36703
rect 28684 36672 28733 36700
rect 28684 36660 28690 36672
rect 28721 36669 28733 36672
rect 28767 36669 28779 36703
rect 28721 36663 28779 36669
rect 28994 36660 29000 36712
rect 29052 36700 29058 36712
rect 29181 36703 29239 36709
rect 29181 36700 29193 36703
rect 29052 36672 29193 36700
rect 29052 36660 29058 36672
rect 29181 36669 29193 36672
rect 29227 36669 29239 36703
rect 29181 36663 29239 36669
rect 29270 36660 29276 36712
rect 29328 36700 29334 36712
rect 29641 36703 29699 36709
rect 29641 36700 29653 36703
rect 29328 36672 29653 36700
rect 29328 36660 29334 36672
rect 29641 36669 29653 36672
rect 29687 36669 29699 36703
rect 34330 36700 34336 36712
rect 34291 36672 34336 36700
rect 29641 36663 29699 36669
rect 34330 36660 34336 36672
rect 34388 36660 34394 36712
rect 34425 36703 34483 36709
rect 34425 36669 34437 36703
rect 34471 36700 34483 36703
rect 34790 36700 34796 36712
rect 34471 36672 34796 36700
rect 34471 36669 34483 36672
rect 34425 36663 34483 36669
rect 34790 36660 34796 36672
rect 34848 36660 34854 36712
rect 35176 36700 35204 36808
rect 35802 36796 35808 36808
rect 35860 36796 35866 36848
rect 36354 36836 36360 36848
rect 36315 36808 36360 36836
rect 36354 36796 36360 36808
rect 36412 36836 36418 36848
rect 37461 36839 37519 36845
rect 37461 36836 37473 36839
rect 36412 36808 37473 36836
rect 36412 36796 36418 36808
rect 37461 36805 37473 36808
rect 37507 36805 37519 36839
rect 37461 36799 37519 36805
rect 37553 36839 37611 36845
rect 37553 36805 37565 36839
rect 37599 36836 37611 36839
rect 37734 36836 37740 36848
rect 37599 36808 37740 36836
rect 37599 36805 37611 36808
rect 37553 36799 37611 36805
rect 37734 36796 37740 36808
rect 37792 36836 37798 36848
rect 40402 36836 40408 36848
rect 37792 36808 40408 36836
rect 37792 36796 37798 36808
rect 40402 36796 40408 36808
rect 40460 36796 40466 36848
rect 40586 36796 40592 36848
rect 40644 36836 40650 36848
rect 41138 36836 41144 36848
rect 40644 36808 41144 36836
rect 40644 36796 40650 36808
rect 41138 36796 41144 36808
rect 41196 36796 41202 36848
rect 41414 36796 41420 36848
rect 41472 36836 41478 36848
rect 41472 36808 44588 36836
rect 41472 36796 41478 36808
rect 35250 36728 35256 36780
rect 35308 36768 35314 36780
rect 35618 36768 35624 36780
rect 35308 36740 35624 36768
rect 35308 36728 35314 36740
rect 35618 36728 35624 36740
rect 35676 36728 35682 36780
rect 36170 36768 36176 36780
rect 36131 36740 36176 36768
rect 36170 36728 36176 36740
rect 36228 36728 36234 36780
rect 36446 36768 36452 36780
rect 36407 36740 36452 36768
rect 36446 36728 36452 36740
rect 36504 36728 36510 36780
rect 36538 36728 36544 36780
rect 36596 36768 36602 36780
rect 37277 36771 37335 36777
rect 36596 36740 36641 36768
rect 36596 36728 36602 36740
rect 37277 36737 37289 36771
rect 37323 36737 37335 36771
rect 37277 36731 37335 36737
rect 35345 36703 35403 36709
rect 35345 36700 35357 36703
rect 35176 36672 35357 36700
rect 35345 36669 35357 36672
rect 35391 36669 35403 36703
rect 35345 36663 35403 36669
rect 35437 36703 35495 36709
rect 35437 36669 35449 36703
rect 35483 36669 35495 36703
rect 35437 36663 35495 36669
rect 35529 36703 35587 36709
rect 35529 36669 35541 36703
rect 35575 36700 35587 36703
rect 35710 36700 35716 36712
rect 35575 36672 35716 36700
rect 35575 36669 35587 36672
rect 35529 36663 35587 36669
rect 31297 36635 31355 36641
rect 26620 36604 28396 36632
rect 28460 36604 30788 36632
rect 26620 36576 26648 36604
rect 25130 36524 25136 36576
rect 25188 36564 25194 36576
rect 25777 36567 25835 36573
rect 25777 36564 25789 36567
rect 25188 36536 25789 36564
rect 25188 36524 25194 36536
rect 25777 36533 25789 36536
rect 25823 36533 25835 36567
rect 25777 36527 25835 36533
rect 26145 36567 26203 36573
rect 26145 36533 26157 36567
rect 26191 36564 26203 36567
rect 26602 36564 26608 36576
rect 26191 36536 26608 36564
rect 26191 36533 26203 36536
rect 26145 36527 26203 36533
rect 26602 36524 26608 36536
rect 26660 36524 26666 36576
rect 27798 36524 27804 36576
rect 27856 36564 27862 36576
rect 28261 36567 28319 36573
rect 28261 36564 28273 36567
rect 27856 36536 28273 36564
rect 27856 36524 27862 36536
rect 28261 36533 28273 36536
rect 28307 36533 28319 36567
rect 28368 36564 28396 36604
rect 28629 36567 28687 36573
rect 28629 36564 28641 36567
rect 28368 36536 28641 36564
rect 28261 36527 28319 36533
rect 28629 36533 28641 36536
rect 28675 36564 28687 36567
rect 29549 36567 29607 36573
rect 29549 36564 29561 36567
rect 28675 36536 29561 36564
rect 28675 36533 28687 36536
rect 28629 36527 28687 36533
rect 29549 36533 29561 36536
rect 29595 36564 29607 36567
rect 29822 36564 29828 36576
rect 29595 36536 29828 36564
rect 29595 36533 29607 36536
rect 29549 36527 29607 36533
rect 29822 36524 29828 36536
rect 29880 36524 29886 36576
rect 30466 36524 30472 36576
rect 30524 36564 30530 36576
rect 30650 36564 30656 36576
rect 30524 36536 30656 36564
rect 30524 36524 30530 36536
rect 30650 36524 30656 36536
rect 30708 36524 30714 36576
rect 30760 36564 30788 36604
rect 31297 36601 31309 36635
rect 31343 36632 31355 36635
rect 32858 36632 32864 36644
rect 31343 36604 32864 36632
rect 31343 36601 31355 36604
rect 31297 36595 31355 36601
rect 32858 36592 32864 36604
rect 32916 36592 32922 36644
rect 33962 36592 33968 36644
rect 34020 36632 34026 36644
rect 35250 36632 35256 36644
rect 34020 36604 35256 36632
rect 34020 36592 34026 36604
rect 35250 36592 35256 36604
rect 35308 36592 35314 36644
rect 35452 36632 35480 36663
rect 35710 36660 35716 36672
rect 35768 36660 35774 36712
rect 37292 36700 37320 36731
rect 37366 36728 37372 36780
rect 37424 36768 37430 36780
rect 37645 36771 37703 36777
rect 37645 36768 37657 36771
rect 37424 36740 37657 36768
rect 37424 36728 37430 36740
rect 37645 36737 37657 36740
rect 37691 36737 37703 36771
rect 37645 36731 37703 36737
rect 40494 36728 40500 36780
rect 40552 36768 40558 36780
rect 40957 36771 41015 36777
rect 40957 36768 40969 36771
rect 40552 36740 40969 36768
rect 40552 36728 40558 36740
rect 40957 36737 40969 36740
rect 41003 36737 41015 36771
rect 44450 36768 44456 36780
rect 44411 36740 44456 36768
rect 40957 36731 41015 36737
rect 44450 36728 44456 36740
rect 44508 36728 44514 36780
rect 44560 36777 44588 36808
rect 44545 36771 44603 36777
rect 44545 36737 44557 36771
rect 44591 36737 44603 36771
rect 44545 36731 44603 36737
rect 36004 36672 37320 36700
rect 36004 36644 36032 36672
rect 35986 36632 35992 36644
rect 35452 36604 35992 36632
rect 35986 36592 35992 36604
rect 36044 36592 36050 36644
rect 41141 36635 41199 36641
rect 41141 36601 41153 36635
rect 41187 36632 41199 36635
rect 42702 36632 42708 36644
rect 41187 36604 42708 36632
rect 41187 36601 41199 36604
rect 41141 36595 41199 36601
rect 42702 36592 42708 36604
rect 42760 36592 42766 36644
rect 44560 36632 44588 36731
rect 44652 36700 44680 36876
rect 44818 36864 44824 36876
rect 44876 36864 44882 36916
rect 49053 36907 49111 36913
rect 49053 36873 49065 36907
rect 49099 36904 49111 36907
rect 50157 36907 50215 36913
rect 49099 36876 50032 36904
rect 49099 36873 49111 36876
rect 49053 36867 49111 36873
rect 48590 36836 48596 36848
rect 48551 36808 48596 36836
rect 48590 36796 48596 36808
rect 48648 36796 48654 36848
rect 49142 36796 49148 36848
rect 49200 36836 49206 36848
rect 49786 36836 49792 36848
rect 49200 36808 49792 36836
rect 49200 36796 49206 36808
rect 49786 36796 49792 36808
rect 49844 36796 49850 36848
rect 50004 36836 50032 36876
rect 50157 36873 50169 36907
rect 50203 36873 50215 36907
rect 50157 36867 50215 36873
rect 56413 36907 56471 36913
rect 56413 36873 56425 36907
rect 56459 36904 56471 36907
rect 56594 36904 56600 36916
rect 56459 36876 56600 36904
rect 56459 36873 56471 36876
rect 56413 36867 56471 36873
rect 50062 36836 50068 36848
rect 50004 36805 50068 36836
rect 45830 36728 45836 36780
rect 45888 36768 45894 36780
rect 46750 36768 46756 36780
rect 45888 36740 46756 36768
rect 45888 36728 45894 36740
rect 46750 36728 46756 36740
rect 46808 36768 46814 36780
rect 47765 36771 47823 36777
rect 47765 36768 47777 36771
rect 46808 36740 47777 36768
rect 46808 36728 46814 36740
rect 47765 36737 47777 36740
rect 47811 36737 47823 36771
rect 47765 36731 47823 36737
rect 48774 36728 48780 36780
rect 48832 36768 48838 36780
rect 48869 36771 48927 36777
rect 50004 36774 50031 36805
rect 48869 36768 48881 36771
rect 48832 36740 48881 36768
rect 48832 36728 48838 36740
rect 48869 36737 48881 36740
rect 48915 36737 48927 36771
rect 50019 36771 50031 36774
rect 50065 36796 50068 36805
rect 50120 36796 50126 36848
rect 50172 36836 50200 36867
rect 56594 36864 56600 36876
rect 56652 36864 56658 36916
rect 56870 36864 56876 36916
rect 56928 36904 56934 36916
rect 57333 36907 57391 36913
rect 57333 36904 57345 36907
rect 56928 36876 57345 36904
rect 56928 36864 56934 36876
rect 57333 36873 57345 36876
rect 57379 36873 57391 36907
rect 57974 36904 57980 36916
rect 57935 36876 57980 36904
rect 57333 36867 57391 36873
rect 50172 36808 50844 36836
rect 50065 36771 50077 36796
rect 50019 36765 50077 36771
rect 48869 36731 48927 36737
rect 50154 36728 50160 36780
rect 50212 36768 50218 36780
rect 50816 36777 50844 36808
rect 50617 36771 50675 36777
rect 50617 36768 50629 36771
rect 50212 36740 50629 36768
rect 50212 36728 50218 36740
rect 50617 36737 50629 36740
rect 50663 36737 50675 36771
rect 50617 36731 50675 36737
rect 50801 36771 50859 36777
rect 50801 36737 50813 36771
rect 50847 36737 50859 36771
rect 54018 36768 54024 36780
rect 53979 36740 54024 36768
rect 50801 36731 50859 36737
rect 54018 36728 54024 36740
rect 54076 36728 54082 36780
rect 55033 36771 55091 36777
rect 55033 36768 55045 36771
rect 54404 36740 55045 36768
rect 47486 36700 47492 36712
rect 44652 36672 47492 36700
rect 47486 36660 47492 36672
rect 47544 36660 47550 36712
rect 47581 36703 47639 36709
rect 47581 36669 47593 36703
rect 47627 36700 47639 36703
rect 48130 36700 48136 36712
rect 47627 36672 48136 36700
rect 47627 36669 47639 36672
rect 47581 36663 47639 36669
rect 48130 36660 48136 36672
rect 48188 36660 48194 36712
rect 48685 36703 48743 36709
rect 48685 36669 48697 36703
rect 48731 36700 48743 36703
rect 49602 36700 49608 36712
rect 48731 36672 49608 36700
rect 48731 36669 48743 36672
rect 48685 36663 48743 36669
rect 49602 36660 49608 36672
rect 49660 36660 49666 36712
rect 53926 36700 53932 36712
rect 53887 36672 53932 36700
rect 53926 36660 53932 36672
rect 53984 36660 53990 36712
rect 46934 36632 46940 36644
rect 44560 36604 46940 36632
rect 46934 36592 46940 36604
rect 46992 36592 46998 36644
rect 54404 36641 54432 36740
rect 55033 36737 55045 36740
rect 55079 36737 55091 36771
rect 55033 36731 55091 36737
rect 56045 36771 56103 36777
rect 56045 36737 56057 36771
rect 56091 36768 56103 36771
rect 56502 36768 56508 36780
rect 56091 36740 56508 36768
rect 56091 36737 56103 36740
rect 56045 36731 56103 36737
rect 56502 36728 56508 36740
rect 56560 36728 56566 36780
rect 56873 36771 56931 36777
rect 56873 36737 56885 36771
rect 56919 36768 56931 36771
rect 57238 36768 57244 36780
rect 56919 36740 57244 36768
rect 56919 36737 56931 36740
rect 56873 36731 56931 36737
rect 57238 36728 57244 36740
rect 57296 36728 57302 36780
rect 57348 36768 57376 36867
rect 57974 36864 57980 36876
rect 58032 36864 58038 36916
rect 57885 36771 57943 36777
rect 57885 36768 57897 36771
rect 57348 36740 57897 36768
rect 57885 36737 57897 36740
rect 57931 36737 57943 36771
rect 57885 36731 57943 36737
rect 54938 36700 54944 36712
rect 54899 36672 54944 36700
rect 54938 36660 54944 36672
rect 54996 36660 55002 36712
rect 55953 36703 56011 36709
rect 55953 36700 55965 36703
rect 55416 36672 55965 36700
rect 55416 36641 55444 36672
rect 55953 36669 55965 36672
rect 55999 36669 56011 36703
rect 55953 36663 56011 36669
rect 54389 36635 54447 36641
rect 54389 36601 54401 36635
rect 54435 36601 54447 36635
rect 54389 36595 54447 36601
rect 55401 36635 55459 36641
rect 55401 36601 55413 36635
rect 55447 36601 55459 36635
rect 55401 36595 55459 36601
rect 57330 36592 57336 36644
rect 57388 36632 57394 36644
rect 57606 36632 57612 36644
rect 57388 36604 57612 36632
rect 57388 36592 57394 36604
rect 57606 36592 57612 36604
rect 57664 36592 57670 36644
rect 33502 36564 33508 36576
rect 30760 36536 33508 36564
rect 33502 36524 33508 36536
rect 33560 36524 33566 36576
rect 34057 36567 34115 36573
rect 34057 36533 34069 36567
rect 34103 36564 34115 36567
rect 34790 36564 34796 36576
rect 34103 36536 34796 36564
rect 34103 36533 34115 36536
rect 34057 36527 34115 36533
rect 34790 36524 34796 36536
rect 34848 36524 34854 36576
rect 35069 36567 35127 36573
rect 35069 36533 35081 36567
rect 35115 36564 35127 36567
rect 35618 36564 35624 36576
rect 35115 36536 35624 36564
rect 35115 36533 35127 36536
rect 35069 36527 35127 36533
rect 35618 36524 35624 36536
rect 35676 36524 35682 36576
rect 36725 36567 36783 36573
rect 36725 36533 36737 36567
rect 36771 36564 36783 36567
rect 37366 36564 37372 36576
rect 36771 36536 37372 36564
rect 36771 36533 36783 36536
rect 36725 36527 36783 36533
rect 37366 36524 37372 36536
rect 37424 36524 37430 36576
rect 37826 36564 37832 36576
rect 37787 36536 37832 36564
rect 37826 36524 37832 36536
rect 37884 36524 37890 36576
rect 44634 36564 44640 36576
rect 44595 36536 44640 36564
rect 44634 36524 44640 36536
rect 44692 36524 44698 36576
rect 47949 36567 48007 36573
rect 47949 36533 47961 36567
rect 47995 36564 48007 36567
rect 48038 36564 48044 36576
rect 47995 36536 48044 36564
rect 47995 36533 48007 36536
rect 47949 36527 48007 36533
rect 48038 36524 48044 36536
rect 48096 36524 48102 36576
rect 48869 36567 48927 36573
rect 48869 36533 48881 36567
rect 48915 36564 48927 36567
rect 48958 36564 48964 36576
rect 48915 36536 48964 36564
rect 48915 36533 48927 36536
rect 48869 36527 48927 36533
rect 48958 36524 48964 36536
rect 49016 36564 49022 36576
rect 49418 36564 49424 36576
rect 49016 36536 49424 36564
rect 49016 36524 49022 36536
rect 49418 36524 49424 36536
rect 49476 36524 49482 36576
rect 49970 36564 49976 36576
rect 49931 36536 49976 36564
rect 49970 36524 49976 36536
rect 50028 36524 50034 36576
rect 50617 36567 50675 36573
rect 50617 36533 50629 36567
rect 50663 36564 50675 36567
rect 52270 36564 52276 36576
rect 50663 36536 52276 36564
rect 50663 36533 50675 36536
rect 50617 36527 50675 36533
rect 52270 36524 52276 36536
rect 52328 36524 52334 36576
rect 57146 36564 57152 36576
rect 57107 36536 57152 36564
rect 57146 36524 57152 36536
rect 57204 36524 57210 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 26602 36360 26608 36372
rect 26563 36332 26608 36360
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 31570 36360 31576 36372
rect 29564 36332 31576 36360
rect 29564 36233 29592 36332
rect 31570 36320 31576 36332
rect 31628 36320 31634 36372
rect 33965 36363 34023 36369
rect 33965 36329 33977 36363
rect 34011 36360 34023 36363
rect 34146 36360 34152 36372
rect 34011 36332 34152 36360
rect 34011 36329 34023 36332
rect 33965 36323 34023 36329
rect 34146 36320 34152 36332
rect 34204 36320 34210 36372
rect 34514 36320 34520 36372
rect 34572 36360 34578 36372
rect 35710 36360 35716 36372
rect 34572 36332 35113 36360
rect 35671 36332 35716 36360
rect 34572 36320 34578 36332
rect 33870 36252 33876 36304
rect 33928 36292 33934 36304
rect 33928 36264 34928 36292
rect 33928 36252 33934 36264
rect 29549 36227 29607 36233
rect 29549 36193 29561 36227
rect 29595 36193 29607 36227
rect 29822 36224 29828 36236
rect 29783 36196 29828 36224
rect 29549 36187 29607 36193
rect 29822 36184 29828 36196
rect 29880 36184 29886 36236
rect 33045 36227 33103 36233
rect 33045 36224 33057 36227
rect 32692 36196 33057 36224
rect 24397 36159 24455 36165
rect 24397 36125 24409 36159
rect 24443 36156 24455 36159
rect 25038 36156 25044 36168
rect 24443 36128 25044 36156
rect 24443 36125 24455 36128
rect 24397 36119 24455 36125
rect 25038 36116 25044 36128
rect 25096 36116 25102 36168
rect 26421 36159 26479 36165
rect 26421 36125 26433 36159
rect 26467 36125 26479 36159
rect 26421 36119 26479 36125
rect 24664 36091 24722 36097
rect 24664 36057 24676 36091
rect 24710 36088 24722 36091
rect 26050 36088 26056 36100
rect 24710 36060 26056 36088
rect 24710 36057 24722 36060
rect 24664 36051 24722 36057
rect 26050 36048 26056 36060
rect 26108 36048 26114 36100
rect 26436 36088 26464 36119
rect 26694 36116 26700 36168
rect 26752 36156 26758 36168
rect 27522 36156 27528 36168
rect 26752 36128 26797 36156
rect 27483 36128 27528 36156
rect 26752 36116 26758 36128
rect 27522 36116 27528 36128
rect 27580 36116 27586 36168
rect 27798 36165 27804 36168
rect 27792 36156 27804 36165
rect 27759 36128 27804 36156
rect 27792 36119 27804 36128
rect 27798 36116 27804 36119
rect 27856 36116 27862 36168
rect 30929 36159 30987 36165
rect 30929 36125 30941 36159
rect 30975 36156 30987 36159
rect 31018 36156 31024 36168
rect 30975 36128 31024 36156
rect 30975 36125 30987 36128
rect 30929 36119 30987 36125
rect 31018 36116 31024 36128
rect 31076 36156 31082 36168
rect 32692 36156 32720 36196
rect 33045 36193 33057 36196
rect 33091 36224 33103 36227
rect 34698 36224 34704 36236
rect 33091 36196 34704 36224
rect 33091 36193 33103 36196
rect 33045 36187 33103 36193
rect 34698 36184 34704 36196
rect 34756 36184 34762 36236
rect 34900 36233 34928 36264
rect 34974 36252 34980 36304
rect 35032 36252 35038 36304
rect 35085 36292 35113 36332
rect 35710 36320 35716 36332
rect 35768 36320 35774 36372
rect 36446 36320 36452 36372
rect 36504 36360 36510 36372
rect 40310 36360 40316 36372
rect 36504 36332 40316 36360
rect 36504 36320 36510 36332
rect 40310 36320 40316 36332
rect 40368 36320 40374 36372
rect 43438 36360 43444 36372
rect 43399 36332 43444 36360
rect 43438 36320 43444 36332
rect 43496 36320 43502 36372
rect 45554 36360 45560 36372
rect 45515 36332 45560 36360
rect 45554 36320 45560 36332
rect 45612 36320 45618 36372
rect 46017 36363 46075 36369
rect 46017 36329 46029 36363
rect 46063 36360 46075 36363
rect 47581 36363 47639 36369
rect 47581 36360 47593 36363
rect 46063 36332 47593 36360
rect 46063 36329 46075 36332
rect 46017 36323 46075 36329
rect 47581 36329 47593 36332
rect 47627 36329 47639 36363
rect 47581 36323 47639 36329
rect 53653 36363 53711 36369
rect 53653 36329 53665 36363
rect 53699 36360 53711 36363
rect 54938 36360 54944 36372
rect 53699 36332 54944 36360
rect 53699 36329 53711 36332
rect 53653 36323 53711 36329
rect 54938 36320 54944 36332
rect 54996 36320 55002 36372
rect 56410 36360 56416 36372
rect 56371 36332 56416 36360
rect 56410 36320 56416 36332
rect 56468 36320 56474 36372
rect 57238 36360 57244 36372
rect 57199 36332 57244 36360
rect 57238 36320 57244 36332
rect 57296 36320 57302 36372
rect 37274 36292 37280 36304
rect 35085 36264 37280 36292
rect 34885 36227 34943 36233
rect 34885 36193 34897 36227
rect 34931 36193 34943 36227
rect 34885 36187 34943 36193
rect 32858 36156 32864 36168
rect 31076 36128 32720 36156
rect 32819 36128 32864 36156
rect 31076 36116 31082 36128
rect 32858 36116 32864 36128
rect 32916 36116 32922 36168
rect 33962 36156 33968 36168
rect 33923 36128 33968 36156
rect 33962 36116 33968 36128
rect 34020 36116 34026 36168
rect 34149 36159 34207 36165
rect 34149 36125 34161 36159
rect 34195 36125 34207 36159
rect 34149 36119 34207 36125
rect 31196 36091 31254 36097
rect 26436 36060 29040 36088
rect 25498 35980 25504 36032
rect 25556 36020 25562 36032
rect 25777 36023 25835 36029
rect 25777 36020 25789 36023
rect 25556 35992 25789 36020
rect 25556 35980 25562 35992
rect 25777 35989 25789 35992
rect 25823 35989 25835 36023
rect 26234 36020 26240 36032
rect 26195 35992 26240 36020
rect 25777 35983 25835 35989
rect 26234 35980 26240 35992
rect 26292 35980 26298 36032
rect 28626 35980 28632 36032
rect 28684 36020 28690 36032
rect 28905 36023 28963 36029
rect 28905 36020 28917 36023
rect 28684 35992 28917 36020
rect 28684 35980 28690 35992
rect 28905 35989 28917 35992
rect 28951 35989 28963 36023
rect 29012 36020 29040 36060
rect 31196 36057 31208 36091
rect 31242 36088 31254 36091
rect 32122 36088 32128 36100
rect 31242 36060 32128 36088
rect 31242 36057 31254 36060
rect 31196 36051 31254 36057
rect 32122 36048 32128 36060
rect 32180 36048 32186 36100
rect 33226 36088 33232 36100
rect 32232 36060 33232 36088
rect 32232 36020 32260 36060
rect 33226 36048 33232 36060
rect 33284 36048 33290 36100
rect 34164 36088 34192 36119
rect 34514 36116 34520 36168
rect 34572 36156 34578 36168
rect 34790 36156 34796 36168
rect 34572 36128 34796 36156
rect 34572 36116 34578 36128
rect 34790 36116 34796 36128
rect 34848 36116 34854 36168
rect 34983 36165 35011 36252
rect 35085 36233 35113 36264
rect 37274 36252 37280 36264
rect 37332 36252 37338 36304
rect 43993 36295 44051 36301
rect 43993 36292 44005 36295
rect 43272 36264 44005 36292
rect 35069 36227 35127 36233
rect 35069 36193 35081 36227
rect 35115 36193 35127 36227
rect 36078 36224 36084 36236
rect 35069 36187 35127 36193
rect 35728 36196 36084 36224
rect 34977 36159 35035 36165
rect 34977 36125 34989 36159
rect 35023 36125 35035 36159
rect 34977 36119 35035 36125
rect 35161 36159 35219 36165
rect 35161 36125 35173 36159
rect 35207 36125 35219 36159
rect 35161 36119 35219 36125
rect 35176 36088 35204 36119
rect 35250 36116 35256 36168
rect 35308 36156 35314 36168
rect 35728 36165 35756 36196
rect 36078 36184 36084 36196
rect 36136 36184 36142 36236
rect 43272 36233 43300 36264
rect 43993 36261 44005 36264
rect 44039 36261 44051 36295
rect 43993 36255 44051 36261
rect 46845 36295 46903 36301
rect 46845 36261 46857 36295
rect 46891 36261 46903 36295
rect 48317 36295 48375 36301
rect 48317 36292 48329 36295
rect 46845 36255 46903 36261
rect 48148 36264 48329 36292
rect 43257 36227 43315 36233
rect 43257 36193 43269 36227
rect 43303 36193 43315 36227
rect 43257 36187 43315 36193
rect 45925 36227 45983 36233
rect 45925 36193 45937 36227
rect 45971 36224 45983 36227
rect 46860 36224 46888 36255
rect 48038 36224 48044 36236
rect 45971 36196 46796 36224
rect 46860 36196 48044 36224
rect 45971 36193 45983 36196
rect 45925 36187 45983 36193
rect 35713 36159 35771 36165
rect 35713 36156 35725 36159
rect 35308 36128 35725 36156
rect 35308 36116 35314 36128
rect 35713 36125 35725 36128
rect 35759 36125 35771 36159
rect 35713 36119 35771 36125
rect 35897 36159 35955 36165
rect 35897 36125 35909 36159
rect 35943 36156 35955 36159
rect 36814 36156 36820 36168
rect 35943 36128 36820 36156
rect 35943 36125 35955 36128
rect 35897 36119 35955 36125
rect 36814 36116 36820 36128
rect 36872 36116 36878 36168
rect 43162 36156 43168 36168
rect 43123 36128 43168 36156
rect 43162 36116 43168 36128
rect 43220 36116 43226 36168
rect 44266 36156 44272 36168
rect 44227 36128 44272 36156
rect 44266 36116 44272 36128
rect 44324 36116 44330 36168
rect 45278 36116 45284 36168
rect 45336 36156 45342 36168
rect 45833 36159 45891 36165
rect 45833 36156 45845 36159
rect 45336 36128 45845 36156
rect 45336 36116 45342 36128
rect 45833 36125 45845 36128
rect 45879 36125 45891 36159
rect 46106 36156 46112 36168
rect 46067 36128 46112 36156
rect 45833 36119 45891 36125
rect 46106 36116 46112 36128
rect 46164 36116 46170 36168
rect 46198 36116 46204 36168
rect 46256 36156 46262 36168
rect 46293 36159 46351 36165
rect 46293 36156 46305 36159
rect 46256 36128 46305 36156
rect 46256 36116 46262 36128
rect 46293 36125 46305 36128
rect 46339 36125 46351 36159
rect 46768 36156 46796 36196
rect 48038 36184 48044 36196
rect 48096 36184 48102 36236
rect 48148 36156 48176 36264
rect 48317 36261 48329 36264
rect 48363 36261 48375 36295
rect 48317 36255 48375 36261
rect 52733 36295 52791 36301
rect 52733 36261 52745 36295
rect 52779 36292 52791 36295
rect 52779 36264 53328 36292
rect 52779 36261 52791 36264
rect 52733 36255 52791 36261
rect 52270 36224 52276 36236
rect 52231 36196 52276 36224
rect 52270 36184 52276 36196
rect 52328 36184 52334 36236
rect 53300 36233 53328 36264
rect 53285 36227 53343 36233
rect 53285 36193 53297 36227
rect 53331 36193 53343 36227
rect 56134 36224 56140 36236
rect 56095 36196 56140 36224
rect 53285 36187 53343 36193
rect 56134 36184 56140 36196
rect 56192 36184 56198 36236
rect 57054 36184 57060 36236
rect 57112 36184 57118 36236
rect 46768 36128 48176 36156
rect 46293 36119 46351 36125
rect 48222 36116 48228 36168
rect 48280 36156 48286 36168
rect 48593 36159 48651 36165
rect 48280 36128 48325 36156
rect 48280 36116 48286 36128
rect 48593 36125 48605 36159
rect 48639 36125 48651 36159
rect 52362 36156 52368 36168
rect 52323 36128 52368 36156
rect 48593 36119 48651 36125
rect 35986 36088 35992 36100
rect 34164 36060 35112 36088
rect 35176 36060 35992 36088
rect 29012 35992 32260 36020
rect 32309 36023 32367 36029
rect 28905 35983 28963 35989
rect 32309 35989 32321 36023
rect 32355 36020 32367 36023
rect 32398 36020 32404 36032
rect 32355 35992 32404 36020
rect 32355 35989 32367 35992
rect 32309 35983 32367 35989
rect 32398 35980 32404 35992
rect 32456 35980 32462 36032
rect 34701 36023 34759 36029
rect 34701 35989 34713 36023
rect 34747 36020 34759 36023
rect 34790 36020 34796 36032
rect 34747 35992 34796 36020
rect 34747 35989 34759 35992
rect 34701 35983 34759 35989
rect 34790 35980 34796 35992
rect 34848 35980 34854 36032
rect 35084 36020 35112 36060
rect 35986 36048 35992 36060
rect 36044 36048 36050 36100
rect 43993 36091 44051 36097
rect 43993 36057 44005 36091
rect 44039 36088 44051 36091
rect 45462 36088 45468 36100
rect 44039 36060 45468 36088
rect 44039 36057 44051 36060
rect 43993 36051 44051 36057
rect 45462 36048 45468 36060
rect 45520 36048 45526 36100
rect 46845 36091 46903 36097
rect 46845 36057 46857 36091
rect 46891 36088 46903 36091
rect 46934 36088 46940 36100
rect 46891 36060 46940 36088
rect 46891 36057 46903 36060
rect 46845 36051 46903 36057
rect 46934 36048 46940 36060
rect 46992 36048 46998 36100
rect 47305 36091 47363 36097
rect 47305 36057 47317 36091
rect 47351 36088 47363 36091
rect 47670 36088 47676 36100
rect 47351 36060 47676 36088
rect 47351 36057 47363 36060
rect 47305 36051 47363 36057
rect 47670 36048 47676 36060
rect 47728 36088 47734 36100
rect 48608 36088 48636 36119
rect 52362 36116 52368 36128
rect 52420 36116 52426 36168
rect 53377 36159 53435 36165
rect 53377 36125 53389 36159
rect 53423 36125 53435 36159
rect 56042 36156 56048 36168
rect 56003 36128 56048 36156
rect 53377 36119 53435 36125
rect 47728 36060 48636 36088
rect 47728 36048 47734 36060
rect 52086 36048 52092 36100
rect 52144 36088 52150 36100
rect 53392 36088 53420 36119
rect 56042 36116 56048 36128
rect 56100 36116 56106 36168
rect 56873 36159 56931 36165
rect 56873 36125 56885 36159
rect 56919 36156 56931 36159
rect 57072 36156 57100 36184
rect 56919 36128 57100 36156
rect 56919 36125 56931 36128
rect 56873 36119 56931 36125
rect 52144 36060 53420 36088
rect 52144 36048 52150 36060
rect 56962 36048 56968 36100
rect 57020 36088 57026 36100
rect 57057 36091 57115 36097
rect 57057 36088 57069 36091
rect 57020 36060 57069 36088
rect 57020 36048 57026 36060
rect 57057 36057 57069 36060
rect 57103 36057 57115 36091
rect 57057 36051 57115 36057
rect 41690 36020 41696 36032
rect 35084 35992 41696 36020
rect 41690 35980 41696 35992
rect 41748 35980 41754 36032
rect 43530 35980 43536 36032
rect 43588 36020 43594 36032
rect 44177 36023 44235 36029
rect 44177 36020 44189 36023
rect 43588 35992 44189 36020
rect 43588 35980 43594 35992
rect 44177 35989 44189 35992
rect 44223 36020 44235 36023
rect 44450 36020 44456 36032
rect 44223 35992 44456 36020
rect 44223 35989 44235 35992
rect 44177 35983 44235 35989
rect 44450 35980 44456 35992
rect 44508 35980 44514 36032
rect 47397 36023 47455 36029
rect 47397 35989 47409 36023
rect 47443 36020 47455 36023
rect 47486 36020 47492 36032
rect 47443 35992 47492 36020
rect 47443 35989 47455 35992
rect 47397 35983 47455 35989
rect 47486 35980 47492 35992
rect 47544 36020 47550 36032
rect 48501 36023 48559 36029
rect 48501 36020 48513 36023
rect 47544 35992 48513 36020
rect 47544 35980 47550 35992
rect 48501 35989 48513 35992
rect 48547 35989 48559 36023
rect 48501 35983 48559 35989
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 26050 35776 26056 35828
rect 26108 35816 26114 35828
rect 26973 35819 27031 35825
rect 26973 35816 26985 35819
rect 26108 35788 26985 35816
rect 26108 35776 26114 35788
rect 26973 35785 26985 35788
rect 27019 35785 27031 35819
rect 32677 35819 32735 35825
rect 32677 35816 32689 35819
rect 26973 35779 27031 35785
rect 30392 35788 32689 35816
rect 30392 35760 30420 35788
rect 32677 35785 32689 35788
rect 32723 35785 32735 35819
rect 35802 35816 35808 35828
rect 32677 35779 32735 35785
rect 35360 35788 35808 35816
rect 25308 35751 25366 35757
rect 25308 35717 25320 35751
rect 25354 35748 25366 35751
rect 26234 35748 26240 35760
rect 25354 35720 26240 35748
rect 25354 35717 25366 35720
rect 25308 35711 25366 35717
rect 26234 35708 26240 35720
rect 26292 35708 26298 35760
rect 30374 35748 30380 35760
rect 27908 35720 30380 35748
rect 25038 35680 25044 35692
rect 24999 35652 25044 35680
rect 25038 35640 25044 35652
rect 25096 35640 25102 35692
rect 25590 35640 25596 35692
rect 25648 35680 25654 35692
rect 27908 35689 27936 35720
rect 30374 35708 30380 35720
rect 30432 35708 30438 35760
rect 30742 35708 30748 35760
rect 30800 35748 30806 35760
rect 30926 35748 30932 35760
rect 30800 35720 30932 35748
rect 30800 35708 30806 35720
rect 30926 35708 30932 35720
rect 30984 35708 30990 35760
rect 31297 35751 31355 35757
rect 31297 35717 31309 35751
rect 31343 35748 31355 35751
rect 31938 35748 31944 35760
rect 31343 35720 31944 35748
rect 31343 35717 31355 35720
rect 31297 35711 31355 35717
rect 31938 35708 31944 35720
rect 31996 35708 32002 35760
rect 32585 35751 32643 35757
rect 32585 35717 32597 35751
rect 32631 35748 32643 35751
rect 32858 35748 32864 35760
rect 32631 35720 32864 35748
rect 32631 35717 32643 35720
rect 32585 35711 32643 35717
rect 32858 35708 32864 35720
rect 32916 35708 32922 35760
rect 34974 35708 34980 35760
rect 35032 35748 35038 35760
rect 35360 35748 35388 35788
rect 35802 35776 35808 35788
rect 35860 35776 35866 35828
rect 43162 35776 43168 35828
rect 43220 35816 43226 35828
rect 43809 35819 43867 35825
rect 43809 35816 43821 35819
rect 43220 35788 43821 35816
rect 43220 35776 43226 35788
rect 43809 35785 43821 35788
rect 43855 35785 43867 35819
rect 43809 35779 43867 35785
rect 43898 35776 43904 35828
rect 43956 35816 43962 35828
rect 44358 35816 44364 35828
rect 43956 35788 44364 35816
rect 43956 35776 43962 35788
rect 44358 35776 44364 35788
rect 44416 35816 44422 35828
rect 46198 35816 46204 35828
rect 44416 35788 46204 35816
rect 44416 35776 44422 35788
rect 46198 35776 46204 35788
rect 46256 35776 46262 35828
rect 48133 35819 48191 35825
rect 48133 35785 48145 35819
rect 48179 35816 48191 35819
rect 48590 35816 48596 35828
rect 48179 35788 48596 35816
rect 48179 35785 48191 35788
rect 48133 35779 48191 35785
rect 48590 35776 48596 35788
rect 48648 35776 48654 35828
rect 38746 35748 38752 35760
rect 35032 35720 35388 35748
rect 37016 35720 38752 35748
rect 35032 35708 35038 35720
rect 27157 35683 27215 35689
rect 25648 35652 26280 35680
rect 25648 35640 25654 35652
rect 26252 35612 26280 35652
rect 27157 35649 27169 35683
rect 27203 35680 27215 35683
rect 27893 35683 27951 35689
rect 27203 35652 27844 35680
rect 27203 35649 27215 35652
rect 27157 35643 27215 35649
rect 27433 35615 27491 35621
rect 27433 35612 27445 35615
rect 26252 35584 27445 35612
rect 27433 35581 27445 35584
rect 27479 35581 27491 35615
rect 27433 35575 27491 35581
rect 26602 35504 26608 35556
rect 26660 35544 26666 35556
rect 27341 35547 27399 35553
rect 27341 35544 27353 35547
rect 26660 35516 27353 35544
rect 26660 35504 26666 35516
rect 27341 35513 27353 35516
rect 27387 35513 27399 35547
rect 27341 35507 27399 35513
rect 26421 35479 26479 35485
rect 26421 35445 26433 35479
rect 26467 35476 26479 35479
rect 26694 35476 26700 35488
rect 26467 35448 26700 35476
rect 26467 35445 26479 35448
rect 26421 35439 26479 35445
rect 26694 35436 26700 35448
rect 26752 35436 26758 35488
rect 27816 35476 27844 35652
rect 27893 35649 27905 35683
rect 27939 35649 27951 35683
rect 27893 35643 27951 35649
rect 28160 35683 28218 35689
rect 28160 35649 28172 35683
rect 28206 35680 28218 35683
rect 28994 35680 29000 35692
rect 28206 35652 29000 35680
rect 28206 35649 28218 35652
rect 28160 35643 28218 35649
rect 28994 35640 29000 35652
rect 29052 35640 29058 35692
rect 31205 35683 31263 35689
rect 31205 35649 31217 35683
rect 31251 35680 31263 35683
rect 31846 35680 31852 35692
rect 31251 35652 31852 35680
rect 31251 35649 31263 35652
rect 31205 35643 31263 35649
rect 31846 35640 31852 35652
rect 31904 35640 31910 35692
rect 33962 35640 33968 35692
rect 34020 35680 34026 35692
rect 34333 35683 34391 35689
rect 34333 35680 34345 35683
rect 34020 35652 34345 35680
rect 34020 35640 34026 35652
rect 34333 35649 34345 35652
rect 34379 35649 34391 35683
rect 34333 35643 34391 35649
rect 34425 35683 34483 35689
rect 34425 35649 34437 35683
rect 34471 35680 34483 35683
rect 34983 35680 35011 35708
rect 34471 35652 35011 35680
rect 35161 35683 35219 35689
rect 34471 35649 34483 35652
rect 34425 35643 34483 35649
rect 35161 35649 35173 35683
rect 35207 35680 35219 35683
rect 35250 35680 35256 35692
rect 35207 35652 35256 35680
rect 35207 35649 35219 35652
rect 35161 35643 35219 35649
rect 35250 35640 35256 35652
rect 35308 35640 35314 35692
rect 35345 35683 35403 35689
rect 35345 35649 35357 35683
rect 35391 35680 35403 35683
rect 37016 35680 37044 35720
rect 38746 35708 38752 35720
rect 38804 35708 38810 35760
rect 43346 35748 43352 35760
rect 41432 35720 43352 35748
rect 35391 35652 37044 35680
rect 35391 35649 35403 35652
rect 35345 35643 35403 35649
rect 37366 35640 37372 35692
rect 37424 35680 37430 35692
rect 37533 35683 37591 35689
rect 37533 35680 37545 35683
rect 37424 35652 37545 35680
rect 37424 35640 37430 35652
rect 37533 35649 37545 35652
rect 37579 35649 37591 35683
rect 40402 35680 40408 35692
rect 40363 35652 40408 35680
rect 37533 35643 37591 35649
rect 40402 35640 40408 35652
rect 40460 35640 40466 35692
rect 41432 35689 41460 35720
rect 43346 35708 43352 35720
rect 43404 35708 43410 35760
rect 43438 35708 43444 35760
rect 43496 35748 43502 35760
rect 45186 35748 45192 35760
rect 43496 35720 43541 35748
rect 43640 35720 45192 35748
rect 43496 35708 43502 35720
rect 41417 35683 41475 35689
rect 41417 35649 41429 35683
rect 41463 35649 41475 35683
rect 41417 35643 41475 35649
rect 42797 35683 42855 35689
rect 42797 35649 42809 35683
rect 42843 35649 42855 35683
rect 42797 35643 42855 35649
rect 42981 35683 43039 35689
rect 42981 35649 42993 35683
rect 43027 35680 43039 35683
rect 43530 35680 43536 35692
rect 43027 35652 43536 35680
rect 43027 35649 43039 35652
rect 42981 35643 43039 35649
rect 31478 35612 31484 35624
rect 31439 35584 31484 35612
rect 31478 35572 31484 35584
rect 31536 35572 31542 35624
rect 32950 35572 32956 35624
rect 33008 35612 33014 35624
rect 34517 35615 34575 35621
rect 34517 35612 34529 35615
rect 33008 35584 34529 35612
rect 33008 35572 33014 35584
rect 34517 35581 34529 35584
rect 34563 35581 34575 35615
rect 34517 35575 34575 35581
rect 34609 35615 34667 35621
rect 34609 35581 34621 35615
rect 34655 35612 34667 35615
rect 35526 35612 35532 35624
rect 34655 35584 35532 35612
rect 34655 35581 34667 35584
rect 34609 35575 34667 35581
rect 33042 35544 33048 35556
rect 28828 35516 33048 35544
rect 28828 35476 28856 35516
rect 33042 35504 33048 35516
rect 33100 35504 33106 35556
rect 34532 35544 34560 35575
rect 35526 35572 35532 35584
rect 35584 35572 35590 35624
rect 37274 35612 37280 35624
rect 37235 35584 37280 35612
rect 37274 35572 37280 35584
rect 37332 35572 37338 35624
rect 40497 35615 40555 35621
rect 40497 35581 40509 35615
rect 40543 35612 40555 35615
rect 41506 35612 41512 35624
rect 40543 35584 41512 35612
rect 40543 35581 40555 35584
rect 40497 35575 40555 35581
rect 41506 35572 41512 35584
rect 41564 35572 41570 35624
rect 41690 35612 41696 35624
rect 41651 35584 41696 35612
rect 41690 35572 41696 35584
rect 41748 35572 41754 35624
rect 42812 35612 42840 35643
rect 43530 35640 43536 35652
rect 43588 35640 43594 35692
rect 43640 35689 43668 35720
rect 45186 35708 45192 35720
rect 45244 35708 45250 35760
rect 45281 35751 45339 35757
rect 45281 35717 45293 35751
rect 45327 35748 45339 35751
rect 46290 35748 46296 35760
rect 45327 35720 46296 35748
rect 45327 35717 45339 35720
rect 45281 35711 45339 35717
rect 46290 35708 46296 35720
rect 46348 35708 46354 35760
rect 49326 35708 49332 35760
rect 49384 35748 49390 35760
rect 49789 35751 49847 35757
rect 49789 35748 49801 35751
rect 49384 35720 49801 35748
rect 49384 35708 49390 35720
rect 49789 35717 49801 35720
rect 49835 35717 49847 35751
rect 49789 35711 49847 35717
rect 49878 35708 49884 35760
rect 49936 35748 49942 35760
rect 49989 35751 50047 35757
rect 49989 35748 50001 35751
rect 49936 35720 50001 35748
rect 49936 35708 49942 35720
rect 49989 35717 50001 35720
rect 50035 35717 50047 35751
rect 49989 35711 50047 35717
rect 51166 35708 51172 35760
rect 51224 35748 51230 35760
rect 51629 35751 51687 35757
rect 51629 35748 51641 35751
rect 51224 35720 51641 35748
rect 51224 35708 51230 35720
rect 51629 35717 51641 35720
rect 51675 35717 51687 35751
rect 51629 35711 51687 35717
rect 55217 35751 55275 35757
rect 55217 35717 55229 35751
rect 55263 35748 55275 35751
rect 56778 35748 56784 35760
rect 55263 35720 56784 35748
rect 55263 35717 55275 35720
rect 55217 35711 55275 35717
rect 56778 35708 56784 35720
rect 56836 35708 56842 35760
rect 43625 35683 43683 35689
rect 43625 35649 43637 35683
rect 43671 35649 43683 35683
rect 43625 35643 43683 35649
rect 44082 35640 44088 35692
rect 44140 35680 44146 35692
rect 44266 35680 44272 35692
rect 44140 35652 44272 35680
rect 44140 35640 44146 35652
rect 44266 35640 44272 35652
rect 44324 35640 44330 35692
rect 44450 35680 44456 35692
rect 44411 35652 44456 35680
rect 44450 35640 44456 35652
rect 44508 35640 44514 35692
rect 45002 35640 45008 35692
rect 45060 35680 45066 35692
rect 45097 35683 45155 35689
rect 45097 35680 45109 35683
rect 45060 35652 45109 35680
rect 45060 35640 45066 35652
rect 45097 35649 45109 35652
rect 45143 35649 45155 35683
rect 45097 35643 45155 35649
rect 45373 35683 45431 35689
rect 45373 35649 45385 35683
rect 45419 35680 45431 35683
rect 46382 35680 46388 35692
rect 45419 35652 46388 35680
rect 45419 35649 45431 35652
rect 45373 35643 45431 35649
rect 46382 35640 46388 35652
rect 46440 35640 46446 35692
rect 48041 35683 48099 35689
rect 48041 35649 48053 35683
rect 48087 35680 48099 35683
rect 48406 35680 48412 35692
rect 48087 35652 48412 35680
rect 48087 35649 48099 35652
rect 48041 35643 48099 35649
rect 48406 35640 48412 35652
rect 48464 35640 48470 35692
rect 49234 35640 49240 35692
rect 49292 35680 49298 35692
rect 50706 35680 50712 35692
rect 49292 35652 50712 35680
rect 49292 35640 49298 35652
rect 50706 35640 50712 35652
rect 50764 35640 50770 35692
rect 51442 35680 51448 35692
rect 51403 35652 51448 35680
rect 51442 35640 51448 35652
rect 51500 35640 51506 35692
rect 51721 35683 51779 35689
rect 51721 35649 51733 35683
rect 51767 35649 51779 35683
rect 51721 35643 51779 35649
rect 55401 35683 55459 35689
rect 55401 35649 55413 35683
rect 55447 35649 55459 35683
rect 56134 35680 56140 35692
rect 56095 35652 56140 35680
rect 55401 35643 55459 35649
rect 44100 35612 44128 35640
rect 42812 35584 44128 35612
rect 44358 35572 44364 35624
rect 44416 35612 44422 35624
rect 46106 35612 46112 35624
rect 44416 35584 46112 35612
rect 44416 35572 44422 35584
rect 46106 35572 46112 35584
rect 46164 35572 46170 35624
rect 48424 35612 48452 35640
rect 48590 35612 48596 35624
rect 48424 35584 48596 35612
rect 48590 35572 48596 35584
rect 48648 35572 48654 35624
rect 51626 35572 51632 35624
rect 51684 35612 51690 35624
rect 51736 35612 51764 35643
rect 51684 35584 51764 35612
rect 51684 35572 51690 35584
rect 36170 35544 36176 35556
rect 34532 35516 36176 35544
rect 36170 35504 36176 35516
rect 36228 35504 36234 35556
rect 41233 35547 41291 35553
rect 41233 35513 41245 35547
rect 41279 35544 41291 35547
rect 55416 35544 55444 35643
rect 56134 35640 56140 35652
rect 56192 35640 56198 35692
rect 41279 35516 55444 35544
rect 41279 35513 41291 35516
rect 41233 35507 41291 35513
rect 29270 35476 29276 35488
rect 27816 35448 28856 35476
rect 29231 35448 29276 35476
rect 29270 35436 29276 35448
rect 29328 35436 29334 35488
rect 30837 35479 30895 35485
rect 30837 35445 30849 35479
rect 30883 35476 30895 35479
rect 33226 35476 33232 35488
rect 30883 35448 33232 35476
rect 30883 35445 30895 35448
rect 30837 35439 30895 35445
rect 33226 35436 33232 35448
rect 33284 35436 33290 35488
rect 34146 35476 34152 35488
rect 34107 35448 34152 35476
rect 34146 35436 34152 35448
rect 34204 35436 34210 35488
rect 35161 35479 35219 35485
rect 35161 35445 35173 35479
rect 35207 35476 35219 35479
rect 35986 35476 35992 35488
rect 35207 35448 35992 35476
rect 35207 35445 35219 35448
rect 35161 35439 35219 35445
rect 35986 35436 35992 35448
rect 36044 35436 36050 35488
rect 38657 35479 38715 35485
rect 38657 35445 38669 35479
rect 38703 35476 38715 35479
rect 38746 35476 38752 35488
rect 38703 35448 38752 35476
rect 38703 35445 38715 35448
rect 38657 35439 38715 35445
rect 38746 35436 38752 35448
rect 38804 35436 38810 35488
rect 40681 35479 40739 35485
rect 40681 35445 40693 35479
rect 40727 35476 40739 35479
rect 40954 35476 40960 35488
rect 40727 35448 40960 35476
rect 40727 35445 40739 35448
rect 40681 35439 40739 35445
rect 40954 35436 40960 35448
rect 41012 35436 41018 35488
rect 41322 35436 41328 35488
rect 41380 35476 41386 35488
rect 41601 35479 41659 35485
rect 41601 35476 41613 35479
rect 41380 35448 41613 35476
rect 41380 35436 41386 35448
rect 41601 35445 41613 35448
rect 41647 35445 41659 35479
rect 42886 35476 42892 35488
rect 42847 35448 42892 35476
rect 41601 35439 41659 35445
rect 42886 35436 42892 35448
rect 42944 35436 42950 35488
rect 43622 35436 43628 35488
rect 43680 35476 43686 35488
rect 44637 35479 44695 35485
rect 44637 35476 44649 35479
rect 43680 35448 44649 35476
rect 43680 35436 43686 35448
rect 44637 35445 44649 35448
rect 44683 35445 44695 35479
rect 45094 35476 45100 35488
rect 45055 35448 45100 35476
rect 44637 35439 44695 35445
rect 45094 35436 45100 35448
rect 45152 35436 45158 35488
rect 49050 35436 49056 35488
rect 49108 35476 49114 35488
rect 49973 35479 50031 35485
rect 49973 35476 49985 35479
rect 49108 35448 49985 35476
rect 49108 35436 49114 35448
rect 49973 35445 49985 35448
rect 50019 35445 50031 35479
rect 50154 35476 50160 35488
rect 50115 35448 50160 35476
rect 49973 35439 50031 35445
rect 50154 35436 50160 35448
rect 50212 35436 50218 35488
rect 50614 35436 50620 35488
rect 50672 35476 50678 35488
rect 50801 35479 50859 35485
rect 50801 35476 50813 35479
rect 50672 35448 50813 35476
rect 50672 35436 50678 35448
rect 50801 35445 50813 35448
rect 50847 35445 50859 35479
rect 50801 35439 50859 35445
rect 51445 35479 51503 35485
rect 51445 35445 51457 35479
rect 51491 35476 51503 35479
rect 53374 35476 53380 35488
rect 51491 35448 53380 35476
rect 51491 35445 51503 35448
rect 51445 35439 51503 35445
rect 53374 35436 53380 35448
rect 53432 35436 53438 35488
rect 55585 35479 55643 35485
rect 55585 35445 55597 35479
rect 55631 35476 55643 35479
rect 56042 35476 56048 35488
rect 55631 35448 56048 35476
rect 55631 35445 55643 35448
rect 55585 35439 55643 35445
rect 56042 35436 56048 35448
rect 56100 35476 56106 35488
rect 56229 35479 56287 35485
rect 56229 35476 56241 35479
rect 56100 35448 56241 35476
rect 56100 35436 56106 35448
rect 56229 35445 56241 35448
rect 56275 35445 56287 35479
rect 56229 35439 56287 35445
rect 56318 35436 56324 35488
rect 56376 35476 56382 35488
rect 56597 35479 56655 35485
rect 56597 35476 56609 35479
rect 56376 35448 56609 35476
rect 56376 35436 56382 35448
rect 56597 35445 56609 35448
rect 56643 35445 56655 35479
rect 56597 35439 56655 35445
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 25038 35272 25044 35284
rect 24872 35244 25044 35272
rect 24872 35145 24900 35244
rect 25038 35232 25044 35244
rect 25096 35272 25102 35284
rect 27341 35275 27399 35281
rect 27341 35272 27353 35275
rect 25096 35244 27353 35272
rect 25096 35232 25102 35244
rect 27341 35241 27353 35244
rect 27387 35272 27399 35275
rect 27522 35272 27528 35284
rect 27387 35244 27528 35272
rect 27387 35241 27399 35244
rect 27341 35235 27399 35241
rect 27522 35232 27528 35244
rect 27580 35232 27586 35284
rect 30006 35232 30012 35284
rect 30064 35272 30070 35284
rect 32401 35275 32459 35281
rect 32401 35272 32413 35275
rect 30064 35244 32413 35272
rect 30064 35232 30070 35244
rect 32401 35241 32413 35244
rect 32447 35272 32459 35275
rect 32582 35272 32588 35284
rect 32447 35244 32588 35272
rect 32447 35241 32459 35244
rect 32401 35235 32459 35241
rect 32582 35232 32588 35244
rect 32640 35232 32646 35284
rect 40497 35275 40555 35281
rect 40497 35241 40509 35275
rect 40543 35272 40555 35275
rect 41046 35272 41052 35284
rect 40543 35244 41052 35272
rect 40543 35241 40555 35244
rect 40497 35235 40555 35241
rect 41046 35232 41052 35244
rect 41104 35232 41110 35284
rect 41874 35272 41880 35284
rect 41835 35244 41880 35272
rect 41874 35232 41880 35244
rect 41932 35272 41938 35284
rect 42702 35272 42708 35284
rect 41932 35244 42708 35272
rect 41932 35232 41938 35244
rect 42702 35232 42708 35244
rect 42760 35232 42766 35284
rect 47210 35272 47216 35284
rect 42812 35244 47072 35272
rect 47171 35244 47216 35272
rect 26237 35207 26295 35213
rect 26237 35173 26249 35207
rect 26283 35204 26295 35207
rect 26326 35204 26332 35216
rect 26283 35176 26332 35204
rect 26283 35173 26295 35176
rect 26237 35167 26295 35173
rect 26326 35164 26332 35176
rect 26384 35164 26390 35216
rect 29825 35207 29883 35213
rect 29825 35173 29837 35207
rect 29871 35204 29883 35207
rect 30926 35204 30932 35216
rect 29871 35176 30932 35204
rect 29871 35173 29883 35176
rect 29825 35167 29883 35173
rect 30926 35164 30932 35176
rect 30984 35164 30990 35216
rect 42812 35204 42840 35244
rect 42628 35176 42840 35204
rect 24857 35139 24915 35145
rect 24857 35105 24869 35139
rect 24903 35105 24915 35139
rect 28166 35136 28172 35148
rect 28127 35108 28172 35136
rect 24857 35099 24915 35105
rect 28166 35096 28172 35108
rect 28224 35096 28230 35148
rect 30469 35139 30527 35145
rect 30469 35105 30481 35139
rect 30515 35136 30527 35139
rect 30742 35136 30748 35148
rect 30515 35108 30748 35136
rect 30515 35105 30527 35108
rect 30469 35099 30527 35105
rect 30742 35096 30748 35108
rect 30800 35096 30806 35148
rect 31018 35136 31024 35148
rect 30979 35108 31024 35136
rect 31018 35096 31024 35108
rect 31076 35096 31082 35148
rect 34698 35136 34704 35148
rect 34659 35108 34704 35136
rect 34698 35096 34704 35108
rect 34756 35096 34762 35148
rect 40954 35136 40960 35148
rect 40915 35108 40960 35136
rect 40954 35096 40960 35108
rect 41012 35096 41018 35148
rect 41046 35096 41052 35148
rect 41104 35136 41110 35148
rect 42518 35136 42524 35148
rect 41104 35108 42524 35136
rect 41104 35096 41110 35108
rect 42518 35096 42524 35108
rect 42576 35096 42582 35148
rect 25130 35077 25136 35080
rect 25124 35068 25136 35077
rect 25091 35040 25136 35068
rect 25124 35031 25136 35040
rect 25130 35028 25136 35031
rect 25188 35028 25194 35080
rect 27246 35068 27252 35080
rect 27207 35040 27252 35068
rect 27246 35028 27252 35040
rect 27304 35028 27310 35080
rect 27614 35028 27620 35080
rect 27672 35068 27678 35080
rect 28445 35071 28503 35077
rect 28445 35068 28457 35071
rect 27672 35040 28457 35068
rect 27672 35028 27678 35040
rect 28445 35037 28457 35040
rect 28491 35037 28503 35071
rect 28445 35031 28503 35037
rect 30285 35071 30343 35077
rect 30285 35037 30297 35071
rect 30331 35068 30343 35071
rect 30834 35068 30840 35080
rect 30331 35040 30840 35068
rect 30331 35037 30343 35040
rect 30285 35031 30343 35037
rect 30834 35028 30840 35040
rect 30892 35028 30898 35080
rect 34716 35068 34744 35096
rect 37185 35071 37243 35077
rect 37185 35068 37197 35071
rect 34716 35040 37197 35068
rect 37185 35037 37197 35040
rect 37231 35068 37243 35071
rect 37274 35068 37280 35080
rect 37231 35040 37280 35068
rect 37231 35037 37243 35040
rect 37185 35031 37243 35037
rect 37274 35028 37280 35040
rect 37332 35028 37338 35080
rect 37452 35071 37510 35077
rect 37452 35037 37464 35071
rect 37498 35068 37510 35071
rect 37826 35068 37832 35080
rect 37498 35040 37832 35068
rect 37498 35037 37510 35040
rect 37452 35031 37510 35037
rect 37826 35028 37832 35040
rect 37884 35028 37890 35080
rect 38654 35028 38660 35080
rect 38712 35068 38718 35080
rect 38712 35040 41276 35068
rect 38712 35028 38718 35040
rect 31288 35003 31346 35009
rect 31288 34969 31300 35003
rect 31334 35000 31346 35003
rect 31938 35000 31944 35012
rect 31334 34972 31944 35000
rect 31334 34969 31346 34972
rect 31288 34963 31346 34969
rect 31938 34960 31944 34972
rect 31996 34960 32002 35012
rect 34968 35003 35026 35009
rect 34968 34969 34980 35003
rect 35014 35000 35026 35003
rect 35434 35000 35440 35012
rect 35014 34972 35440 35000
rect 35014 34969 35026 34972
rect 34968 34963 35026 34969
rect 35434 34960 35440 34972
rect 35492 34960 35498 35012
rect 40865 35003 40923 35009
rect 40865 34969 40877 35003
rect 40911 35000 40923 35003
rect 41248 35000 41276 35040
rect 41322 35028 41328 35080
rect 41380 35068 41386 35080
rect 41693 35071 41751 35077
rect 41693 35068 41705 35071
rect 41380 35040 41705 35068
rect 41380 35028 41386 35040
rect 41693 35037 41705 35040
rect 41739 35037 41751 35071
rect 41693 35031 41751 35037
rect 42628 35000 42656 35176
rect 42886 35164 42892 35216
rect 42944 35204 42950 35216
rect 42944 35176 43760 35204
rect 42944 35164 42950 35176
rect 43073 35139 43131 35145
rect 43073 35105 43085 35139
rect 43119 35136 43131 35139
rect 43346 35136 43352 35148
rect 43119 35108 43352 35136
rect 43119 35105 43131 35108
rect 43073 35099 43131 35105
rect 43346 35096 43352 35108
rect 43404 35096 43410 35148
rect 43622 35136 43628 35148
rect 43583 35108 43628 35136
rect 43622 35096 43628 35108
rect 43680 35096 43686 35148
rect 43732 35145 43760 35176
rect 44008 35176 45232 35204
rect 43717 35139 43775 35145
rect 43717 35105 43729 35139
rect 43763 35105 43775 35139
rect 43717 35099 43775 35105
rect 42705 35071 42763 35077
rect 42705 35037 42717 35071
rect 42751 35068 42763 35071
rect 42981 35071 43039 35077
rect 42751 35040 42932 35068
rect 42751 35037 42763 35040
rect 42705 35031 42763 35037
rect 40911 34972 41184 35000
rect 41248 34972 42656 35000
rect 42904 35000 42932 35040
rect 42981 35037 42993 35071
rect 43027 35068 43039 35071
rect 44008 35068 44036 35176
rect 44361 35139 44419 35145
rect 44361 35105 44373 35139
rect 44407 35136 44419 35139
rect 45094 35136 45100 35148
rect 44407 35108 45100 35136
rect 44407 35105 44419 35108
rect 44361 35099 44419 35105
rect 45094 35096 45100 35108
rect 45152 35096 45158 35148
rect 45204 35136 45232 35176
rect 45462 35164 45468 35216
rect 45520 35204 45526 35216
rect 46109 35207 46167 35213
rect 46109 35204 46121 35207
rect 45520 35176 46121 35204
rect 45520 35164 45526 35176
rect 46109 35173 46121 35176
rect 46155 35173 46167 35207
rect 47044 35204 47072 35244
rect 47210 35232 47216 35244
rect 47268 35232 47274 35284
rect 49050 35232 49056 35284
rect 49108 35272 49114 35284
rect 49237 35275 49295 35281
rect 49237 35272 49249 35275
rect 49108 35244 49249 35272
rect 49108 35232 49114 35244
rect 49237 35241 49249 35244
rect 49283 35241 49295 35275
rect 49237 35235 49295 35241
rect 50709 35275 50767 35281
rect 50709 35241 50721 35275
rect 50755 35272 50767 35275
rect 52086 35272 52092 35284
rect 50755 35244 52092 35272
rect 50755 35241 50767 35244
rect 50709 35235 50767 35241
rect 52086 35232 52092 35244
rect 52144 35232 52150 35284
rect 52181 35275 52239 35281
rect 52181 35241 52193 35275
rect 52227 35272 52239 35275
rect 52362 35272 52368 35284
rect 52227 35244 52368 35272
rect 52227 35241 52239 35244
rect 52181 35235 52239 35241
rect 52362 35232 52368 35244
rect 52420 35232 52426 35284
rect 57146 35232 57152 35284
rect 57204 35272 57210 35284
rect 57241 35275 57299 35281
rect 57241 35272 57253 35275
rect 57204 35244 57253 35272
rect 57204 35232 57210 35244
rect 57241 35241 57253 35244
rect 57287 35241 57299 35275
rect 57241 35235 57299 35241
rect 48682 35204 48688 35216
rect 47044 35176 48688 35204
rect 46109 35167 46167 35173
rect 48682 35164 48688 35176
rect 48740 35164 48746 35216
rect 51166 35204 51172 35216
rect 51046 35176 51172 35204
rect 51046 35136 51074 35176
rect 51166 35164 51172 35176
rect 51224 35204 51230 35216
rect 52270 35204 52276 35216
rect 51224 35176 52276 35204
rect 51224 35164 51230 35176
rect 52270 35164 52276 35176
rect 52328 35164 52334 35216
rect 51258 35136 51264 35148
rect 45204 35108 51074 35136
rect 51219 35108 51264 35136
rect 51258 35096 51264 35108
rect 51316 35096 51322 35148
rect 52546 35136 52552 35148
rect 52507 35108 52552 35136
rect 52546 35096 52552 35108
rect 52604 35096 52610 35148
rect 43027 35040 44036 35068
rect 44085 35071 44143 35077
rect 43027 35037 43039 35040
rect 42981 35031 43039 35037
rect 44085 35037 44097 35071
rect 44131 35068 44143 35071
rect 44266 35068 44272 35080
rect 44131 35040 44272 35068
rect 44131 35037 44143 35040
rect 44085 35031 44143 35037
rect 44266 35028 44272 35040
rect 44324 35068 44330 35080
rect 45002 35068 45008 35080
rect 44324 35040 45008 35068
rect 44324 35028 44330 35040
rect 45002 35028 45008 35040
rect 45060 35028 45066 35080
rect 45649 35071 45707 35077
rect 45649 35068 45661 35071
rect 45112 35040 45661 35068
rect 43254 35000 43260 35012
rect 42904 34972 43260 35000
rect 40911 34969 40923 34972
rect 40865 34963 40923 34969
rect 30098 34892 30104 34944
rect 30156 34932 30162 34944
rect 30193 34935 30251 34941
rect 30193 34932 30205 34935
rect 30156 34904 30205 34932
rect 30156 34892 30162 34904
rect 30193 34901 30205 34904
rect 30239 34901 30251 34935
rect 30193 34895 30251 34901
rect 36081 34935 36139 34941
rect 36081 34901 36093 34935
rect 36127 34932 36139 34935
rect 37182 34932 37188 34944
rect 36127 34904 37188 34932
rect 36127 34901 36139 34904
rect 36081 34895 36139 34901
rect 37182 34892 37188 34904
rect 37240 34892 37246 34944
rect 38565 34935 38623 34941
rect 38565 34901 38577 34935
rect 38611 34932 38623 34935
rect 39114 34932 39120 34944
rect 38611 34904 39120 34932
rect 38611 34901 38623 34904
rect 38565 34895 38623 34901
rect 39114 34892 39120 34904
rect 39172 34892 39178 34944
rect 41156 34932 41184 34972
rect 43254 34960 43260 34972
rect 43312 34960 43318 35012
rect 43714 34960 43720 35012
rect 43772 35000 43778 35012
rect 44177 35003 44235 35009
rect 44177 35000 44189 35003
rect 43772 34972 44189 35000
rect 43772 34960 43778 34972
rect 44177 34969 44189 34972
rect 44223 34969 44235 35003
rect 44177 34963 44235 34969
rect 44910 34960 44916 35012
rect 44968 35000 44974 35012
rect 45112 35000 45140 35040
rect 45649 35037 45661 35040
rect 45695 35068 45707 35071
rect 45695 35040 46336 35068
rect 45695 35037 45707 35040
rect 45649 35031 45707 35037
rect 44968 34972 45140 35000
rect 45465 35003 45523 35009
rect 44968 34960 44974 34972
rect 45465 34969 45477 35003
rect 45511 34969 45523 35003
rect 45465 34963 45523 34969
rect 41414 34932 41420 34944
rect 41156 34904 41420 34932
rect 41414 34892 41420 34904
rect 41472 34892 41478 34944
rect 43272 34932 43300 34960
rect 45480 34932 45508 34963
rect 45922 34960 45928 35012
rect 45980 35000 45986 35012
rect 46109 35003 46167 35009
rect 46109 35000 46121 35003
rect 45980 34972 46121 35000
rect 45980 34960 45986 34972
rect 46109 34969 46121 34972
rect 46155 34969 46167 35003
rect 46308 35000 46336 35040
rect 46382 35028 46388 35080
rect 46440 35068 46446 35080
rect 47121 35071 47179 35077
rect 46440 35040 46485 35068
rect 46440 35028 46446 35040
rect 47121 35037 47133 35071
rect 47167 35037 47179 35071
rect 47121 35031 47179 35037
rect 47136 35000 47164 35031
rect 47210 35028 47216 35080
rect 47268 35068 47274 35080
rect 47305 35071 47363 35077
rect 47305 35068 47317 35071
rect 47268 35040 47317 35068
rect 47268 35028 47274 35040
rect 47305 35037 47317 35040
rect 47351 35037 47363 35071
rect 49970 35068 49976 35080
rect 47305 35031 47363 35037
rect 49160 35040 49976 35068
rect 47394 35000 47400 35012
rect 46308 34972 46428 35000
rect 47136 34972 47400 35000
rect 46109 34963 46167 34969
rect 46290 34932 46296 34944
rect 43272 34904 45508 34932
rect 46251 34904 46296 34932
rect 46290 34892 46296 34904
rect 46348 34892 46354 34944
rect 46400 34932 46428 34972
rect 47394 34960 47400 34972
rect 47452 34960 47458 35012
rect 48958 34960 48964 35012
rect 49016 35000 49022 35012
rect 49160 35009 49188 35040
rect 49970 35028 49976 35040
rect 50028 35028 50034 35080
rect 50154 35028 50160 35080
rect 50212 35068 50218 35080
rect 51077 35071 51135 35077
rect 51077 35068 51089 35071
rect 50212 35040 51089 35068
rect 50212 35028 50218 35040
rect 51077 35037 51089 35040
rect 51123 35037 51135 35071
rect 51077 35031 51135 35037
rect 52365 35071 52423 35077
rect 52365 35037 52377 35071
rect 52411 35037 52423 35071
rect 52365 35031 52423 35037
rect 49145 35003 49203 35009
rect 49145 35000 49157 35003
rect 49016 34972 49157 35000
rect 49016 34960 49022 34972
rect 49145 34969 49157 34972
rect 49191 34969 49203 35003
rect 52380 35000 52408 35031
rect 52454 35028 52460 35080
rect 52512 35068 52518 35080
rect 52512 35040 52557 35068
rect 52512 35028 52518 35040
rect 52638 35028 52644 35080
rect 52696 35068 52702 35080
rect 53193 35071 53251 35077
rect 53193 35068 53205 35071
rect 52696 35040 53205 35068
rect 52696 35028 52702 35040
rect 53193 35037 53205 35040
rect 53239 35037 53251 35071
rect 53374 35068 53380 35080
rect 53335 35040 53380 35068
rect 53193 35031 53251 35037
rect 53374 35028 53380 35040
rect 53432 35028 53438 35080
rect 56229 35071 56287 35077
rect 56229 35037 56241 35071
rect 56275 35068 56287 35071
rect 56318 35068 56324 35080
rect 56275 35040 56324 35068
rect 56275 35037 56287 35040
rect 56229 35031 56287 35037
rect 56318 35028 56324 35040
rect 56376 35028 56382 35080
rect 56413 35071 56471 35077
rect 56413 35037 56425 35071
rect 56459 35037 56471 35071
rect 56962 35068 56968 35080
rect 56923 35040 56968 35068
rect 56413 35031 56471 35037
rect 49145 34963 49203 34969
rect 49252 34972 51856 35000
rect 52380 34972 53328 35000
rect 49252 34932 49280 34972
rect 51166 34932 51172 34944
rect 46400 34904 49280 34932
rect 51127 34904 51172 34932
rect 51166 34892 51172 34904
rect 51224 34892 51230 34944
rect 51828 34932 51856 34972
rect 52454 34932 52460 34944
rect 51828 34904 52460 34932
rect 52454 34892 52460 34904
rect 52512 34932 52518 34944
rect 52730 34932 52736 34944
rect 52512 34904 52736 34932
rect 52512 34892 52518 34904
rect 52730 34892 52736 34904
rect 52788 34892 52794 34944
rect 53300 34941 53328 34972
rect 55582 34960 55588 35012
rect 55640 35000 55646 35012
rect 56428 35000 56456 35031
rect 56962 35028 56968 35040
rect 57020 35028 57026 35080
rect 57054 35028 57060 35080
rect 57112 35068 57118 35080
rect 57112 35040 57157 35068
rect 57112 35028 57118 35040
rect 55640 34972 56456 35000
rect 55640 34960 55646 34972
rect 53285 34935 53343 34941
rect 53285 34901 53297 34935
rect 53331 34932 53343 34935
rect 53466 34932 53472 34944
rect 53331 34904 53472 34932
rect 53331 34901 53343 34904
rect 53285 34895 53343 34901
rect 53466 34892 53472 34904
rect 53524 34892 53530 34944
rect 56413 34935 56471 34941
rect 56413 34901 56425 34935
rect 56459 34932 56471 34935
rect 56980 34932 57008 35028
rect 56459 34904 57008 34932
rect 56459 34901 56471 34904
rect 56413 34895 56471 34901
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 31573 34731 31631 34737
rect 31573 34697 31585 34731
rect 31619 34728 31631 34731
rect 31846 34728 31852 34740
rect 31619 34700 31852 34728
rect 31619 34697 31631 34700
rect 31573 34691 31631 34697
rect 31846 34688 31852 34700
rect 31904 34688 31910 34740
rect 38654 34728 38660 34740
rect 38615 34700 38660 34728
rect 38654 34688 38660 34700
rect 38712 34688 38718 34740
rect 40402 34688 40408 34740
rect 40460 34728 40466 34740
rect 41049 34731 41107 34737
rect 41049 34728 41061 34731
rect 40460 34700 41061 34728
rect 40460 34688 40466 34700
rect 41049 34697 41061 34700
rect 41095 34728 41107 34731
rect 41095 34700 41460 34728
rect 41095 34697 41107 34700
rect 41049 34691 41107 34697
rect 30374 34620 30380 34672
rect 30432 34660 30438 34672
rect 35710 34660 35716 34672
rect 30432 34632 35716 34660
rect 30432 34620 30438 34632
rect 28166 34592 28172 34604
rect 28127 34564 28172 34592
rect 28166 34552 28172 34564
rect 28224 34552 28230 34604
rect 30193 34595 30251 34601
rect 30193 34561 30205 34595
rect 30239 34592 30251 34595
rect 30392 34592 30420 34620
rect 30239 34564 30420 34592
rect 30460 34595 30518 34601
rect 30239 34561 30251 34564
rect 30193 34555 30251 34561
rect 30460 34561 30472 34595
rect 30506 34592 30518 34595
rect 30506 34564 31432 34592
rect 30506 34561 30518 34564
rect 30460 34555 30518 34561
rect 27614 34484 27620 34536
rect 27672 34524 27678 34536
rect 27985 34527 28043 34533
rect 27985 34524 27997 34527
rect 27672 34496 27997 34524
rect 27672 34484 27678 34496
rect 27985 34493 27997 34496
rect 28031 34493 28043 34527
rect 27985 34487 28043 34493
rect 27706 34348 27712 34400
rect 27764 34388 27770 34400
rect 28353 34391 28411 34397
rect 28353 34388 28365 34391
rect 27764 34360 28365 34388
rect 27764 34348 27770 34360
rect 28353 34357 28365 34360
rect 28399 34357 28411 34391
rect 31404 34388 31432 34564
rect 32306 34552 32312 34604
rect 32364 34592 32370 34604
rect 32582 34592 32588 34604
rect 32364 34564 32409 34592
rect 32543 34564 32588 34592
rect 32364 34552 32370 34564
rect 32582 34552 32588 34564
rect 32640 34552 32646 34604
rect 33226 34592 33232 34604
rect 33187 34564 33232 34592
rect 33226 34552 33232 34564
rect 33284 34552 33290 34604
rect 34072 34601 34100 34632
rect 35710 34620 35716 34632
rect 35768 34660 35774 34672
rect 37544 34663 37602 34669
rect 35768 34632 37320 34660
rect 35768 34620 35774 34632
rect 34057 34595 34115 34601
rect 34057 34561 34069 34595
rect 34103 34561 34115 34595
rect 34057 34555 34115 34561
rect 34146 34552 34152 34604
rect 34204 34592 34210 34604
rect 37292 34601 37320 34632
rect 37544 34629 37556 34663
rect 37590 34660 37602 34663
rect 38378 34660 38384 34672
rect 37590 34632 38384 34660
rect 37590 34629 37602 34632
rect 37544 34623 37602 34629
rect 38378 34620 38384 34632
rect 38436 34620 38442 34672
rect 40310 34620 40316 34672
rect 40368 34660 40374 34672
rect 41322 34660 41328 34672
rect 40368 34632 41328 34660
rect 40368 34620 40374 34632
rect 41322 34620 41328 34632
rect 41380 34620 41386 34672
rect 41432 34660 41460 34700
rect 41506 34688 41512 34740
rect 41564 34728 41570 34740
rect 42981 34731 43039 34737
rect 42981 34728 42993 34731
rect 41564 34700 42993 34728
rect 41564 34688 41570 34700
rect 42981 34697 42993 34700
rect 43027 34697 43039 34731
rect 42981 34691 43039 34697
rect 43349 34731 43407 34737
rect 43349 34697 43361 34731
rect 43395 34728 43407 34731
rect 44358 34728 44364 34740
rect 43395 34700 43944 34728
rect 44319 34700 44364 34728
rect 43395 34697 43407 34700
rect 43349 34691 43407 34697
rect 41693 34663 41751 34669
rect 41693 34660 41705 34663
rect 41432 34632 41705 34660
rect 41693 34629 41705 34632
rect 41739 34660 41751 34663
rect 42794 34660 42800 34672
rect 41739 34632 42800 34660
rect 41739 34629 41751 34632
rect 41693 34623 41751 34629
rect 42794 34620 42800 34632
rect 42852 34620 42858 34672
rect 42886 34620 42892 34672
rect 42944 34660 42950 34672
rect 43916 34669 43944 34700
rect 44358 34688 44364 34700
rect 44416 34688 44422 34740
rect 44450 34688 44456 34740
rect 44508 34728 44514 34740
rect 46477 34731 46535 34737
rect 46477 34728 46489 34731
rect 44508 34700 46489 34728
rect 44508 34688 44514 34700
rect 46477 34697 46489 34700
rect 46523 34697 46535 34731
rect 46477 34691 46535 34697
rect 49053 34731 49111 34737
rect 49053 34697 49065 34731
rect 49099 34728 49111 34731
rect 49878 34728 49884 34740
rect 49099 34700 49884 34728
rect 49099 34697 49111 34700
rect 49053 34691 49111 34697
rect 49878 34688 49884 34700
rect 49936 34688 49942 34740
rect 49970 34688 49976 34740
rect 50028 34728 50034 34740
rect 50028 34700 50384 34728
rect 50028 34688 50034 34700
rect 43901 34663 43959 34669
rect 42944 34632 43484 34660
rect 42944 34620 42950 34632
rect 34313 34595 34371 34601
rect 34313 34592 34325 34595
rect 34204 34564 34325 34592
rect 34204 34552 34210 34564
rect 34313 34561 34325 34564
rect 34359 34561 34371 34595
rect 34313 34555 34371 34561
rect 37277 34595 37335 34601
rect 37277 34561 37289 34595
rect 37323 34561 37335 34595
rect 40402 34592 40408 34604
rect 37277 34555 37335 34561
rect 37384 34564 38332 34592
rect 40363 34564 40408 34592
rect 31478 34484 31484 34536
rect 31536 34524 31542 34536
rect 32493 34527 32551 34533
rect 32493 34524 32505 34527
rect 31536 34496 32505 34524
rect 31536 34484 31542 34496
rect 32493 34493 32505 34496
rect 32539 34493 32551 34527
rect 35526 34524 35532 34536
rect 32493 34487 32551 34493
rect 35452 34496 35532 34524
rect 31938 34416 31944 34468
rect 31996 34456 32002 34468
rect 35452 34465 35480 34496
rect 35526 34484 35532 34496
rect 35584 34524 35590 34536
rect 37384 34524 37412 34564
rect 35584 34496 37412 34524
rect 38304 34524 38332 34564
rect 40402 34552 40408 34564
rect 40460 34552 40466 34604
rect 40681 34595 40739 34601
rect 40681 34561 40693 34595
rect 40727 34592 40739 34595
rect 41414 34592 41420 34604
rect 40727 34564 41420 34592
rect 40727 34561 40739 34564
rect 40681 34555 40739 34561
rect 41414 34552 41420 34564
rect 41472 34552 41478 34604
rect 41506 34552 41512 34604
rect 41564 34592 41570 34604
rect 43165 34595 43223 34601
rect 41564 34564 41609 34592
rect 41564 34552 41570 34564
rect 43165 34561 43177 34595
rect 43211 34592 43223 34595
rect 43346 34592 43352 34604
rect 43211 34564 43352 34592
rect 43211 34561 43223 34564
rect 43165 34555 43223 34561
rect 43346 34552 43352 34564
rect 43404 34552 43410 34604
rect 43456 34601 43484 34632
rect 43901 34629 43913 34663
rect 43947 34660 43959 34663
rect 45925 34663 45983 34669
rect 45925 34660 45937 34663
rect 43947 34632 45937 34660
rect 43947 34629 43959 34632
rect 43901 34623 43959 34629
rect 45925 34629 45937 34632
rect 45971 34629 45983 34663
rect 47486 34660 47492 34672
rect 45925 34623 45983 34629
rect 46676 34632 47492 34660
rect 43441 34595 43499 34601
rect 43441 34561 43453 34595
rect 43487 34561 43499 34595
rect 44174 34592 44180 34604
rect 44135 34564 44180 34592
rect 43441 34555 43499 34561
rect 44174 34552 44180 34564
rect 44232 34552 44238 34604
rect 44450 34552 44456 34604
rect 44508 34592 44514 34604
rect 44913 34595 44971 34601
rect 44913 34592 44925 34595
rect 44508 34564 44925 34592
rect 44508 34552 44514 34564
rect 44913 34561 44925 34564
rect 44959 34592 44971 34595
rect 45094 34592 45100 34604
rect 44959 34564 45100 34592
rect 44959 34561 44971 34564
rect 44913 34555 44971 34561
rect 45094 34552 45100 34564
rect 45152 34552 45158 34604
rect 45186 34552 45192 34604
rect 45244 34592 45250 34604
rect 46676 34601 46704 34632
rect 47486 34620 47492 34632
rect 47544 34620 47550 34672
rect 49789 34663 49847 34669
rect 49789 34660 49801 34663
rect 48884 34632 49801 34660
rect 45833 34595 45891 34601
rect 45244 34564 45289 34592
rect 45244 34552 45250 34564
rect 45833 34561 45845 34595
rect 45879 34561 45891 34595
rect 46017 34595 46075 34601
rect 46017 34592 46029 34595
rect 45833 34555 45891 34561
rect 45940 34564 46029 34592
rect 40494 34524 40500 34536
rect 38304 34496 40500 34524
rect 35584 34484 35590 34496
rect 40494 34484 40500 34496
rect 40552 34484 40558 34536
rect 44085 34527 44143 34533
rect 44085 34524 44097 34527
rect 43640 34496 44097 34524
rect 32125 34459 32183 34465
rect 32125 34456 32137 34459
rect 31996 34428 32137 34456
rect 31996 34416 32002 34428
rect 32125 34425 32137 34428
rect 32171 34425 32183 34459
rect 32125 34419 32183 34425
rect 35437 34459 35495 34465
rect 35437 34425 35449 34459
rect 35483 34425 35495 34459
rect 35437 34419 35495 34425
rect 43346 34416 43352 34468
rect 43404 34456 43410 34468
rect 43640 34456 43668 34496
rect 44085 34493 44097 34496
rect 44131 34524 44143 34527
rect 44131 34496 44772 34524
rect 44131 34493 44143 34496
rect 44085 34487 44143 34493
rect 43404 34428 43668 34456
rect 43404 34416 43410 34428
rect 44744 34400 44772 34496
rect 44818 34484 44824 34536
rect 44876 34524 44882 34536
rect 45005 34527 45063 34533
rect 45005 34524 45017 34527
rect 44876 34496 45017 34524
rect 44876 34484 44882 34496
rect 45005 34493 45017 34496
rect 45051 34524 45063 34527
rect 45462 34524 45468 34536
rect 45051 34496 45468 34524
rect 45051 34493 45063 34496
rect 45005 34487 45063 34493
rect 45462 34484 45468 34496
rect 45520 34524 45526 34536
rect 45848 34524 45876 34555
rect 45520 34496 45876 34524
rect 45520 34484 45526 34496
rect 45186 34416 45192 34468
rect 45244 34456 45250 34468
rect 45940 34456 45968 34564
rect 46017 34561 46029 34564
rect 46063 34561 46075 34595
rect 46017 34555 46075 34561
rect 46661 34595 46719 34601
rect 46661 34561 46673 34595
rect 46707 34561 46719 34595
rect 46661 34555 46719 34561
rect 46845 34595 46903 34601
rect 46845 34561 46857 34595
rect 46891 34592 46903 34595
rect 47118 34592 47124 34604
rect 46891 34564 47124 34592
rect 46891 34561 46903 34564
rect 46845 34555 46903 34561
rect 47118 34552 47124 34564
rect 47176 34552 47182 34604
rect 47670 34592 47676 34604
rect 47228 34564 47676 34592
rect 46753 34527 46811 34533
rect 46753 34493 46765 34527
rect 46799 34493 46811 34527
rect 46934 34524 46940 34536
rect 46895 34496 46940 34524
rect 46753 34487 46811 34493
rect 45244 34428 45968 34456
rect 46768 34456 46796 34487
rect 46934 34484 46940 34496
rect 46992 34484 46998 34536
rect 47228 34524 47256 34564
rect 47670 34552 47676 34564
rect 47728 34592 47734 34604
rect 47857 34595 47915 34601
rect 47857 34592 47869 34595
rect 47728 34564 47869 34592
rect 47728 34552 47734 34564
rect 47857 34561 47869 34564
rect 47903 34561 47915 34595
rect 47857 34555 47915 34561
rect 48406 34552 48412 34604
rect 48464 34592 48470 34604
rect 48682 34592 48688 34604
rect 48464 34564 48688 34592
rect 48464 34552 48470 34564
rect 48682 34552 48688 34564
rect 48740 34592 48746 34604
rect 48884 34601 48912 34632
rect 49789 34629 49801 34632
rect 49835 34629 49847 34663
rect 49789 34623 49847 34629
rect 50065 34663 50123 34669
rect 50065 34629 50077 34663
rect 50111 34660 50123 34663
rect 50246 34660 50252 34672
rect 50111 34632 50252 34660
rect 50111 34629 50123 34632
rect 50065 34623 50123 34629
rect 48869 34595 48927 34601
rect 48869 34592 48881 34595
rect 48740 34564 48881 34592
rect 48740 34552 48746 34564
rect 48869 34561 48881 34564
rect 48915 34561 48927 34595
rect 49050 34592 49056 34604
rect 49011 34564 49056 34592
rect 48869 34555 48927 34561
rect 49050 34552 49056 34564
rect 49108 34592 49114 34604
rect 49513 34595 49571 34601
rect 49513 34592 49525 34595
rect 49108 34564 49525 34592
rect 49108 34552 49114 34564
rect 49513 34561 49525 34564
rect 49559 34561 49571 34595
rect 49513 34555 49571 34561
rect 49697 34595 49755 34601
rect 49697 34561 49709 34595
rect 49743 34561 49755 34595
rect 49697 34555 49755 34561
rect 47044 34496 47256 34524
rect 47044 34456 47072 34496
rect 47302 34484 47308 34536
rect 47360 34524 47366 34536
rect 47581 34527 47639 34533
rect 47581 34524 47593 34527
rect 47360 34496 47593 34524
rect 47360 34484 47366 34496
rect 47581 34493 47593 34496
rect 47627 34493 47639 34527
rect 47581 34487 47639 34493
rect 49234 34484 49240 34536
rect 49292 34524 49298 34536
rect 49712 34524 49740 34555
rect 49292 34496 49740 34524
rect 49804 34524 49832 34623
rect 50246 34620 50252 34632
rect 50304 34620 50310 34672
rect 50356 34660 50384 34700
rect 50982 34688 50988 34740
rect 51040 34728 51046 34740
rect 51718 34728 51724 34740
rect 51040 34700 51724 34728
rect 51040 34688 51046 34700
rect 51718 34688 51724 34700
rect 51776 34728 51782 34740
rect 51905 34731 51963 34737
rect 51905 34728 51917 34731
rect 51776 34700 51917 34728
rect 51776 34688 51782 34700
rect 51905 34697 51917 34700
rect 51951 34697 51963 34731
rect 51905 34691 51963 34697
rect 52270 34688 52276 34740
rect 52328 34728 52334 34740
rect 52917 34731 52975 34737
rect 52917 34728 52929 34731
rect 52328 34700 52929 34728
rect 52328 34688 52334 34700
rect 52917 34697 52929 34700
rect 52963 34697 52975 34731
rect 52917 34691 52975 34697
rect 50709 34663 50767 34669
rect 50709 34660 50721 34663
rect 50356 34632 50721 34660
rect 50709 34629 50721 34632
rect 50755 34629 50767 34663
rect 50709 34623 50767 34629
rect 50798 34620 50804 34672
rect 50856 34660 50862 34672
rect 50856 34632 50901 34660
rect 50856 34620 50862 34632
rect 49878 34552 49884 34604
rect 49936 34592 49942 34604
rect 49936 34564 49981 34592
rect 49936 34552 49942 34564
rect 50154 34552 50160 34604
rect 50212 34592 50218 34604
rect 50525 34595 50583 34601
rect 50525 34592 50537 34595
rect 50212 34564 50537 34592
rect 50212 34552 50218 34564
rect 50525 34561 50537 34564
rect 50571 34561 50583 34595
rect 50893 34595 50951 34601
rect 50893 34582 50905 34595
rect 50525 34555 50583 34561
rect 50812 34561 50905 34582
rect 50939 34561 50951 34595
rect 50812 34555 50951 34561
rect 50812 34554 50936 34555
rect 50812 34524 50840 34554
rect 51166 34552 51172 34604
rect 51224 34552 51230 34604
rect 51442 34552 51448 34604
rect 51500 34592 51506 34604
rect 51718 34592 51724 34604
rect 51500 34564 51724 34592
rect 51500 34552 51506 34564
rect 51718 34552 51724 34564
rect 51776 34552 51782 34604
rect 51994 34592 52000 34604
rect 51955 34564 52000 34592
rect 51994 34552 52000 34564
rect 52052 34552 52058 34604
rect 52178 34552 52184 34604
rect 52236 34592 52242 34604
rect 52733 34595 52791 34601
rect 52733 34592 52745 34595
rect 52236 34564 52745 34592
rect 52236 34552 52242 34564
rect 52733 34561 52745 34564
rect 52779 34561 52791 34595
rect 52733 34555 52791 34561
rect 56686 34552 56692 34604
rect 56744 34592 56750 34604
rect 56873 34595 56931 34601
rect 56873 34592 56885 34595
rect 56744 34564 56885 34592
rect 56744 34552 56750 34564
rect 56873 34561 56885 34564
rect 56919 34561 56931 34595
rect 56873 34555 56931 34561
rect 49804 34496 50840 34524
rect 49292 34484 49298 34496
rect 51184 34456 51212 34552
rect 51537 34527 51595 34533
rect 51537 34493 51549 34527
rect 51583 34524 51595 34527
rect 53650 34524 53656 34536
rect 51583 34496 53656 34524
rect 51583 34493 51595 34496
rect 51537 34487 51595 34493
rect 53650 34484 53656 34496
rect 53708 34484 53714 34536
rect 46768 34428 47072 34456
rect 50908 34428 51212 34456
rect 45244 34416 45250 34428
rect 33045 34391 33103 34397
rect 33045 34388 33057 34391
rect 31404 34360 33057 34388
rect 28353 34351 28411 34357
rect 33045 34357 33057 34360
rect 33091 34357 33103 34391
rect 33045 34351 33103 34357
rect 41877 34391 41935 34397
rect 41877 34357 41889 34391
rect 41923 34388 41935 34391
rect 41966 34388 41972 34400
rect 41923 34360 41972 34388
rect 41923 34357 41935 34360
rect 41877 34351 41935 34357
rect 41966 34348 41972 34360
rect 42024 34348 42030 34400
rect 44174 34388 44180 34400
rect 44135 34360 44180 34388
rect 44174 34348 44180 34360
rect 44232 34348 44238 34400
rect 44726 34348 44732 34400
rect 44784 34388 44790 34400
rect 44913 34391 44971 34397
rect 44913 34388 44925 34391
rect 44784 34360 44925 34388
rect 44784 34348 44790 34360
rect 44913 34357 44925 34360
rect 44959 34357 44971 34391
rect 44913 34351 44971 34357
rect 45002 34348 45008 34400
rect 45060 34388 45066 34400
rect 45373 34391 45431 34397
rect 45373 34388 45385 34391
rect 45060 34360 45385 34388
rect 45060 34348 45066 34360
rect 45373 34357 45385 34360
rect 45419 34357 45431 34391
rect 45373 34351 45431 34357
rect 46934 34348 46940 34400
rect 46992 34388 46998 34400
rect 47946 34388 47952 34400
rect 46992 34360 47952 34388
rect 46992 34348 46998 34360
rect 47946 34348 47952 34360
rect 48004 34388 48010 34400
rect 48222 34388 48228 34400
rect 48004 34360 48228 34388
rect 48004 34348 48010 34360
rect 48222 34348 48228 34360
rect 48280 34348 48286 34400
rect 50798 34348 50804 34400
rect 50856 34388 50862 34400
rect 50908 34388 50936 34428
rect 51074 34388 51080 34400
rect 50856 34360 50936 34388
rect 51035 34360 51080 34388
rect 50856 34348 50862 34360
rect 51074 34348 51080 34360
rect 51132 34348 51138 34400
rect 56962 34388 56968 34400
rect 56923 34360 56968 34388
rect 56962 34348 56968 34360
rect 57020 34348 57026 34400
rect 58066 34388 58072 34400
rect 58027 34360 58072 34388
rect 58066 34348 58072 34360
rect 58124 34348 58130 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 28166 34184 28172 34196
rect 28127 34156 28172 34184
rect 28166 34144 28172 34156
rect 28224 34144 28230 34196
rect 39114 34184 39120 34196
rect 39027 34156 39120 34184
rect 39114 34144 39120 34156
rect 39172 34144 39178 34196
rect 40126 34144 40132 34196
rect 40184 34184 40190 34196
rect 40313 34187 40371 34193
rect 40313 34184 40325 34187
rect 40184 34156 40325 34184
rect 40184 34144 40190 34156
rect 40313 34153 40325 34156
rect 40359 34153 40371 34187
rect 43898 34184 43904 34196
rect 40313 34147 40371 34153
rect 41386 34156 43904 34184
rect 39132 34116 39160 34144
rect 41386 34116 41414 34156
rect 43898 34144 43904 34156
rect 43956 34144 43962 34196
rect 44085 34187 44143 34193
rect 44085 34153 44097 34187
rect 44131 34184 44143 34187
rect 45002 34184 45008 34196
rect 44131 34156 45008 34184
rect 44131 34153 44143 34156
rect 44085 34147 44143 34153
rect 45002 34144 45008 34156
rect 45060 34144 45066 34196
rect 45189 34187 45247 34193
rect 45189 34153 45201 34187
rect 45235 34184 45247 34187
rect 46290 34184 46296 34196
rect 45235 34156 46296 34184
rect 45235 34153 45247 34156
rect 45189 34147 45247 34153
rect 46290 34144 46296 34156
rect 46348 34144 46354 34196
rect 47213 34187 47271 34193
rect 47213 34153 47225 34187
rect 47259 34184 47271 34187
rect 47486 34184 47492 34196
rect 47259 34156 47492 34184
rect 47259 34153 47271 34156
rect 47213 34147 47271 34153
rect 47486 34144 47492 34156
rect 47544 34144 47550 34196
rect 47578 34144 47584 34196
rect 47636 34184 47642 34196
rect 51261 34187 51319 34193
rect 47636 34156 51212 34184
rect 47636 34144 47642 34156
rect 43717 34119 43775 34125
rect 39132 34088 41414 34116
rect 41524 34088 42196 34116
rect 25498 34048 25504 34060
rect 25459 34020 25504 34048
rect 25498 34008 25504 34020
rect 25556 34008 25562 34060
rect 25685 34051 25743 34057
rect 25685 34017 25697 34051
rect 25731 34048 25743 34051
rect 28626 34048 28632 34060
rect 25731 34020 26924 34048
rect 28587 34020 28632 34048
rect 25731 34017 25743 34020
rect 25685 34011 25743 34017
rect 26896 33924 26924 34020
rect 28626 34008 28632 34020
rect 28684 34008 28690 34060
rect 28813 34051 28871 34057
rect 28813 34017 28825 34051
rect 28859 34048 28871 34051
rect 30098 34048 30104 34060
rect 28859 34020 30104 34048
rect 28859 34017 28871 34020
rect 28813 34011 28871 34017
rect 27706 33980 27712 33992
rect 27667 33952 27712 33980
rect 27706 33940 27712 33952
rect 27764 33940 27770 33992
rect 25409 33915 25467 33921
rect 25409 33881 25421 33915
rect 25455 33912 25467 33915
rect 26050 33912 26056 33924
rect 25455 33884 26056 33912
rect 25455 33881 25467 33884
rect 25409 33875 25467 33881
rect 26050 33872 26056 33884
rect 26108 33872 26114 33924
rect 26878 33872 26884 33924
rect 26936 33912 26942 33924
rect 28828 33912 28856 34011
rect 30098 34008 30104 34020
rect 30156 34008 30162 34060
rect 30374 34008 30380 34060
rect 30432 34048 30438 34060
rect 30745 34051 30803 34057
rect 30745 34048 30757 34051
rect 30432 34020 30757 34048
rect 30432 34008 30438 34020
rect 30745 34017 30757 34020
rect 30791 34017 30803 34051
rect 34698 34048 34704 34060
rect 34659 34020 34704 34048
rect 30745 34011 30803 34017
rect 34698 34008 34704 34020
rect 34756 34008 34762 34060
rect 38654 34008 38660 34060
rect 38712 34048 38718 34060
rect 39025 34051 39083 34057
rect 39025 34048 39037 34051
rect 38712 34020 39037 34048
rect 38712 34008 38718 34020
rect 39025 34017 39037 34020
rect 39071 34017 39083 34051
rect 39025 34011 39083 34017
rect 40957 34051 41015 34057
rect 40957 34017 40969 34051
rect 41003 34048 41015 34051
rect 41046 34048 41052 34060
rect 41003 34020 41052 34048
rect 41003 34017 41015 34020
rect 40957 34011 41015 34017
rect 41046 34008 41052 34020
rect 41104 34008 41110 34060
rect 41524 34057 41552 34088
rect 41509 34051 41567 34057
rect 41509 34017 41521 34051
rect 41555 34048 41567 34051
rect 41598 34048 41604 34060
rect 41555 34020 41604 34048
rect 41555 34017 41567 34020
rect 41509 34011 41567 34017
rect 41598 34008 41604 34020
rect 41656 34008 41662 34060
rect 41966 34048 41972 34060
rect 41927 34020 41972 34048
rect 41966 34008 41972 34020
rect 42024 34008 42030 34060
rect 42168 34048 42196 34088
rect 43717 34085 43729 34119
rect 43763 34116 43775 34119
rect 43806 34116 43812 34128
rect 43763 34088 43812 34116
rect 43763 34085 43775 34088
rect 43717 34079 43775 34085
rect 43806 34076 43812 34088
rect 43864 34076 43870 34128
rect 44266 34116 44272 34128
rect 44227 34088 44272 34116
rect 44266 34076 44272 34088
rect 44324 34076 44330 34128
rect 45373 34119 45431 34125
rect 45373 34085 45385 34119
rect 45419 34085 45431 34119
rect 45373 34079 45431 34085
rect 44174 34048 44180 34060
rect 42168 34020 44180 34048
rect 44174 34008 44180 34020
rect 44232 34008 44238 34060
rect 34606 33940 34612 33992
rect 34664 33980 34670 33992
rect 34957 33983 35015 33989
rect 34957 33980 34969 33983
rect 34664 33952 34969 33980
rect 34664 33940 34670 33952
rect 34957 33949 34969 33952
rect 35003 33949 35015 33983
rect 34957 33943 35015 33949
rect 38746 33940 38752 33992
rect 38804 33980 38810 33992
rect 38933 33983 38991 33989
rect 38933 33980 38945 33983
rect 38804 33952 38945 33980
rect 38804 33940 38810 33952
rect 38933 33949 38945 33952
rect 38979 33980 38991 33983
rect 39114 33980 39120 33992
rect 38979 33952 39120 33980
rect 38979 33949 38991 33952
rect 38933 33943 38991 33949
rect 39114 33940 39120 33952
rect 39172 33940 39178 33992
rect 41874 33980 41880 33992
rect 41835 33952 41880 33980
rect 41874 33940 41880 33952
rect 41932 33940 41938 33992
rect 42978 33940 42984 33992
rect 43036 33980 43042 33992
rect 43993 33983 44051 33989
rect 43993 33980 44005 33983
rect 43036 33952 44005 33980
rect 43036 33940 43042 33952
rect 43993 33949 44005 33952
rect 44039 33949 44051 33983
rect 43993 33943 44051 33949
rect 44453 33983 44511 33989
rect 44453 33949 44465 33983
rect 44499 33980 44511 33983
rect 44910 33980 44916 33992
rect 44499 33952 44916 33980
rect 44499 33949 44511 33952
rect 44453 33943 44511 33949
rect 44910 33940 44916 33952
rect 44968 33940 44974 33992
rect 45094 33940 45100 33992
rect 45152 33980 45158 33992
rect 45388 33980 45416 34079
rect 45738 34076 45744 34128
rect 45796 34116 45802 34128
rect 45796 34088 48636 34116
rect 45796 34076 45802 34088
rect 46934 34008 46940 34060
rect 46992 34048 46998 34060
rect 47210 34048 47216 34060
rect 46992 34020 47216 34048
rect 46992 34008 46998 34020
rect 47210 34008 47216 34020
rect 47268 34048 47274 34060
rect 47489 34051 47547 34057
rect 47489 34048 47501 34051
rect 47268 34020 47501 34048
rect 47268 34008 47274 34020
rect 47489 34017 47501 34020
rect 47535 34017 47547 34051
rect 47489 34011 47547 34017
rect 47673 34051 47731 34057
rect 47673 34017 47685 34051
rect 47719 34048 47731 34051
rect 48314 34048 48320 34060
rect 47719 34020 48320 34048
rect 47719 34017 47731 34020
rect 47673 34011 47731 34017
rect 48314 34008 48320 34020
rect 48372 34008 48378 34060
rect 45152 33952 45416 33980
rect 45152 33940 45158 33952
rect 46474 33940 46480 33992
rect 46532 33980 46538 33992
rect 46753 33983 46811 33989
rect 46532 33952 46577 33980
rect 46532 33940 46538 33952
rect 46753 33949 46765 33983
rect 46799 33980 46811 33983
rect 47394 33980 47400 33992
rect 46799 33952 47400 33980
rect 46799 33949 46811 33952
rect 46753 33943 46811 33949
rect 47394 33940 47400 33952
rect 47452 33940 47458 33992
rect 47581 33983 47639 33989
rect 47581 33949 47593 33983
rect 47627 33980 47639 33983
rect 47854 33980 47860 33992
rect 47627 33952 47860 33980
rect 47627 33949 47639 33952
rect 47581 33943 47639 33949
rect 26936 33884 28856 33912
rect 26936 33872 26942 33884
rect 30742 33872 30748 33924
rect 30800 33912 30806 33924
rect 30990 33915 31048 33921
rect 30990 33912 31002 33915
rect 30800 33884 31002 33912
rect 30800 33872 30806 33884
rect 30990 33881 31002 33884
rect 31036 33881 31048 33915
rect 30990 33875 31048 33881
rect 40773 33915 40831 33921
rect 40773 33881 40785 33915
rect 40819 33912 40831 33915
rect 42153 33915 42211 33921
rect 42153 33912 42165 33915
rect 40819 33884 42165 33912
rect 40819 33881 40831 33884
rect 40773 33875 40831 33881
rect 42153 33881 42165 33884
rect 42199 33881 42211 33915
rect 42153 33875 42211 33881
rect 42518 33872 42524 33924
rect 42576 33912 42582 33924
rect 42705 33915 42763 33921
rect 42705 33912 42717 33915
rect 42576 33884 42717 33912
rect 42576 33872 42582 33884
rect 42705 33881 42717 33884
rect 42751 33881 42763 33915
rect 45002 33912 45008 33924
rect 44963 33884 45008 33912
rect 42705 33875 42763 33881
rect 45002 33872 45008 33884
rect 45060 33872 45066 33924
rect 45221 33915 45279 33921
rect 45221 33881 45233 33915
rect 45267 33912 45279 33915
rect 45370 33912 45376 33924
rect 45267 33884 45376 33912
rect 45267 33881 45279 33884
rect 45221 33875 45279 33881
rect 45370 33872 45376 33884
rect 45428 33872 45434 33924
rect 46293 33915 46351 33921
rect 46293 33881 46305 33915
rect 46339 33912 46351 33915
rect 47302 33912 47308 33924
rect 46339 33884 47308 33912
rect 46339 33881 46351 33884
rect 46293 33875 46351 33881
rect 47302 33872 47308 33884
rect 47360 33872 47366 33924
rect 24118 33804 24124 33856
rect 24176 33844 24182 33856
rect 25041 33847 25099 33853
rect 25041 33844 25053 33847
rect 24176 33816 25053 33844
rect 24176 33804 24182 33816
rect 25041 33813 25053 33816
rect 25087 33813 25099 33847
rect 27522 33844 27528 33856
rect 27483 33816 27528 33844
rect 25041 33807 25099 33813
rect 27522 33804 27528 33816
rect 27580 33804 27586 33856
rect 28537 33847 28595 33853
rect 28537 33813 28549 33847
rect 28583 33844 28595 33847
rect 29086 33844 29092 33856
rect 28583 33816 29092 33844
rect 28583 33813 28595 33816
rect 28537 33807 28595 33813
rect 29086 33804 29092 33816
rect 29144 33804 29150 33856
rect 29914 33804 29920 33856
rect 29972 33844 29978 33856
rect 32125 33847 32183 33853
rect 32125 33844 32137 33847
rect 29972 33816 32137 33844
rect 29972 33804 29978 33816
rect 32125 33813 32137 33816
rect 32171 33813 32183 33847
rect 36078 33844 36084 33856
rect 36039 33816 36084 33844
rect 32125 33807 32183 33813
rect 36078 33804 36084 33816
rect 36136 33804 36142 33856
rect 39298 33844 39304 33856
rect 39259 33816 39304 33844
rect 39298 33804 39304 33816
rect 39356 33804 39362 33856
rect 40678 33844 40684 33856
rect 40639 33816 40684 33844
rect 40678 33804 40684 33816
rect 40736 33804 40742 33856
rect 40862 33804 40868 33856
rect 40920 33844 40926 33856
rect 41230 33844 41236 33856
rect 40920 33816 41236 33844
rect 40920 33804 40926 33816
rect 41230 33804 41236 33816
rect 41288 33844 41294 33856
rect 42794 33844 42800 33856
rect 41288 33816 42800 33844
rect 41288 33804 41294 33816
rect 42794 33804 42800 33816
rect 42852 33804 42858 33856
rect 46661 33847 46719 33853
rect 46661 33813 46673 33847
rect 46707 33844 46719 33847
rect 46934 33844 46940 33856
rect 46707 33816 46940 33844
rect 46707 33813 46719 33816
rect 46661 33807 46719 33813
rect 46934 33804 46940 33816
rect 46992 33804 46998 33856
rect 47210 33804 47216 33856
rect 47268 33844 47274 33856
rect 47596 33844 47624 33943
rect 47854 33940 47860 33952
rect 47912 33940 47918 33992
rect 48406 33980 48412 33992
rect 48367 33952 48412 33980
rect 48406 33940 48412 33952
rect 48464 33940 48470 33992
rect 47268 33816 47624 33844
rect 47268 33804 47274 33816
rect 48406 33804 48412 33856
rect 48464 33844 48470 33856
rect 48501 33847 48559 33853
rect 48501 33844 48513 33847
rect 48464 33816 48513 33844
rect 48464 33804 48470 33816
rect 48501 33813 48513 33816
rect 48547 33813 48559 33847
rect 48608 33844 48636 34088
rect 51184 34048 51212 34156
rect 51261 34153 51273 34187
rect 51307 34184 51319 34187
rect 51350 34184 51356 34196
rect 51307 34156 51356 34184
rect 51307 34153 51319 34156
rect 51261 34147 51319 34153
rect 51350 34144 51356 34156
rect 51408 34144 51414 34196
rect 51626 34144 51632 34196
rect 51684 34184 51690 34196
rect 51997 34187 52055 34193
rect 51997 34184 52009 34187
rect 51684 34156 52009 34184
rect 51684 34144 51690 34156
rect 51997 34153 52009 34156
rect 52043 34153 52055 34187
rect 51997 34147 52055 34153
rect 52181 34187 52239 34193
rect 52181 34153 52193 34187
rect 52227 34184 52239 34187
rect 52638 34184 52644 34196
rect 52227 34156 52644 34184
rect 52227 34153 52239 34156
rect 52181 34147 52239 34153
rect 52638 34144 52644 34156
rect 52696 34144 52702 34196
rect 54478 34184 54484 34196
rect 54439 34156 54484 34184
rect 54478 34144 54484 34156
rect 54536 34144 54542 34196
rect 55861 34187 55919 34193
rect 55861 34153 55873 34187
rect 55907 34184 55919 34187
rect 56134 34184 56140 34196
rect 55907 34156 56140 34184
rect 55907 34153 55919 34156
rect 55861 34147 55919 34153
rect 56134 34144 56140 34156
rect 56192 34144 56198 34196
rect 58066 34116 58072 34128
rect 56336 34088 58072 34116
rect 51626 34048 51632 34060
rect 51184 34020 51632 34048
rect 51626 34008 51632 34020
rect 51684 34008 51690 34060
rect 52546 34008 52552 34060
rect 52604 34048 52610 34060
rect 52730 34048 52736 34060
rect 52604 34020 52736 34048
rect 52604 34008 52610 34020
rect 52730 34008 52736 34020
rect 52788 34048 52794 34060
rect 53466 34048 53472 34060
rect 52788 34020 52868 34048
rect 53427 34020 53472 34048
rect 52788 34008 52794 34020
rect 49878 33980 49884 33992
rect 49344 33952 49884 33980
rect 49344 33924 49372 33952
rect 49878 33940 49884 33952
rect 49936 33940 49942 33992
rect 50062 33940 50068 33992
rect 50120 33980 50126 33992
rect 50120 33952 50292 33980
rect 50120 33940 50126 33952
rect 49326 33912 49332 33924
rect 49287 33884 49332 33912
rect 49326 33872 49332 33884
rect 49384 33872 49390 33924
rect 49513 33915 49571 33921
rect 49513 33881 49525 33915
rect 49559 33912 49571 33915
rect 50154 33912 50160 33924
rect 49559 33884 50160 33912
rect 49559 33881 49571 33884
rect 49513 33875 49571 33881
rect 50154 33872 50160 33884
rect 50212 33872 50218 33924
rect 50264 33912 50292 33952
rect 50890 33940 50896 33992
rect 50948 33980 50954 33992
rect 52362 33980 52368 33992
rect 50948 33952 52368 33980
rect 50948 33940 50954 33952
rect 52362 33940 52368 33952
rect 52420 33940 52426 33992
rect 52454 33940 52460 33992
rect 52512 33980 52518 33992
rect 52840 33989 52868 34020
rect 53466 34008 53472 34020
rect 53524 34008 53530 34060
rect 56336 34057 56364 34088
rect 58066 34076 58072 34088
rect 58124 34076 58130 34128
rect 56321 34051 56379 34057
rect 56321 34017 56333 34051
rect 56367 34017 56379 34051
rect 56321 34011 56379 34017
rect 56505 34051 56563 34057
rect 56505 34017 56517 34051
rect 56551 34048 56563 34051
rect 56962 34048 56968 34060
rect 56551 34020 56968 34048
rect 56551 34017 56563 34020
rect 56505 34011 56563 34017
rect 56962 34008 56968 34020
rect 57020 34008 57026 34060
rect 57882 34048 57888 34060
rect 57843 34020 57888 34048
rect 57882 34008 57888 34020
rect 57940 34008 57946 34060
rect 52641 33983 52699 33989
rect 52641 33980 52653 33983
rect 52512 33952 52653 33980
rect 52512 33940 52518 33952
rect 52641 33949 52653 33952
rect 52687 33949 52699 33983
rect 52641 33943 52699 33949
rect 52825 33983 52883 33989
rect 52825 33949 52837 33983
rect 52871 33949 52883 33983
rect 52825 33943 52883 33949
rect 53561 33983 53619 33989
rect 53561 33949 53573 33983
rect 53607 33949 53619 33983
rect 54478 33980 54484 33992
rect 54439 33952 54484 33980
rect 53561 33943 53619 33949
rect 50985 33915 51043 33921
rect 50985 33912 50997 33915
rect 50264 33884 50997 33912
rect 50985 33881 50997 33884
rect 51031 33881 51043 33915
rect 50985 33875 51043 33881
rect 51813 33915 51871 33921
rect 51813 33881 51825 33915
rect 51859 33912 51871 33915
rect 52178 33912 52184 33924
rect 51859 33884 52184 33912
rect 51859 33881 51871 33884
rect 51813 33875 51871 33881
rect 52178 33872 52184 33884
rect 52236 33872 52242 33924
rect 52733 33915 52791 33921
rect 52733 33881 52745 33915
rect 52779 33912 52791 33915
rect 53576 33912 53604 33943
rect 54478 33940 54484 33952
rect 54536 33940 54542 33992
rect 54662 33980 54668 33992
rect 54623 33952 54668 33980
rect 54662 33940 54668 33952
rect 54720 33940 54726 33992
rect 55582 33980 55588 33992
rect 55543 33952 55588 33980
rect 55582 33940 55588 33952
rect 55640 33940 55646 33992
rect 55677 33983 55735 33989
rect 55677 33949 55689 33983
rect 55723 33980 55735 33983
rect 55858 33980 55864 33992
rect 55723 33952 55864 33980
rect 55723 33949 55735 33952
rect 55677 33943 55735 33949
rect 55858 33940 55864 33952
rect 55916 33940 55922 33992
rect 52779 33884 53604 33912
rect 52779 33881 52791 33884
rect 52733 33875 52791 33881
rect 51350 33844 51356 33856
rect 48608 33816 51356 33844
rect 48501 33807 48559 33813
rect 51350 33804 51356 33816
rect 51408 33804 51414 33856
rect 51718 33804 51724 33856
rect 51776 33844 51782 33856
rect 52013 33847 52071 33853
rect 52013 33844 52025 33847
rect 51776 33816 52025 33844
rect 51776 33804 51782 33816
rect 52013 33813 52025 33816
rect 52059 33813 52071 33847
rect 52013 33807 52071 33813
rect 53929 33847 53987 33853
rect 53929 33813 53941 33847
rect 53975 33844 53987 33847
rect 55490 33844 55496 33856
rect 53975 33816 55496 33844
rect 53975 33813 53987 33816
rect 53929 33807 53987 33813
rect 55490 33804 55496 33816
rect 55548 33844 55554 33856
rect 56318 33844 56324 33856
rect 55548 33816 56324 33844
rect 55548 33804 55554 33816
rect 56318 33804 56324 33816
rect 56376 33804 56382 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 26053 33643 26111 33649
rect 26053 33609 26065 33643
rect 26099 33640 26111 33643
rect 26326 33640 26332 33652
rect 26099 33612 26332 33640
rect 26099 33609 26111 33612
rect 26053 33603 26111 33609
rect 26326 33600 26332 33612
rect 26384 33600 26390 33652
rect 30742 33640 30748 33652
rect 30703 33612 30748 33640
rect 30742 33600 30748 33612
rect 30800 33600 30806 33652
rect 41598 33640 41604 33652
rect 41559 33612 41604 33640
rect 41598 33600 41604 33612
rect 41656 33600 41662 33652
rect 42794 33600 42800 33652
rect 42852 33600 42858 33652
rect 42978 33640 42984 33652
rect 42939 33612 42984 33640
rect 42978 33600 42984 33612
rect 43036 33600 43042 33652
rect 44269 33643 44327 33649
rect 44269 33609 44281 33643
rect 44315 33640 44327 33643
rect 45186 33640 45192 33652
rect 44315 33612 45192 33640
rect 44315 33609 44327 33612
rect 44269 33603 44327 33609
rect 45186 33600 45192 33612
rect 45244 33600 45250 33652
rect 45554 33640 45560 33652
rect 45515 33612 45560 33640
rect 45554 33600 45560 33612
rect 45612 33600 45618 33652
rect 46474 33600 46480 33652
rect 46532 33640 46538 33652
rect 47210 33640 47216 33652
rect 46532 33612 47216 33640
rect 46532 33600 46538 33612
rect 47210 33600 47216 33612
rect 47268 33600 47274 33652
rect 47302 33600 47308 33652
rect 47360 33640 47366 33652
rect 47673 33643 47731 33649
rect 47673 33640 47685 33643
rect 47360 33612 47685 33640
rect 47360 33600 47366 33612
rect 47673 33609 47685 33612
rect 47719 33609 47731 33643
rect 47673 33603 47731 33609
rect 47857 33643 47915 33649
rect 47857 33609 47869 33643
rect 47903 33609 47915 33643
rect 47857 33603 47915 33609
rect 27522 33532 27528 33584
rect 27580 33572 27586 33584
rect 27770 33575 27828 33581
rect 27770 33572 27782 33575
rect 27580 33544 27782 33572
rect 27580 33532 27586 33544
rect 27770 33541 27782 33544
rect 27816 33541 27828 33575
rect 29914 33572 29920 33584
rect 29875 33544 29920 33572
rect 27770 33535 27828 33541
rect 29914 33532 29920 33544
rect 29972 33532 29978 33584
rect 30098 33572 30104 33584
rect 30059 33544 30104 33572
rect 30098 33532 30104 33544
rect 30156 33532 30162 33584
rect 40957 33575 41015 33581
rect 40957 33541 40969 33575
rect 41003 33572 41015 33575
rect 41322 33572 41328 33584
rect 41003 33544 41328 33572
rect 41003 33541 41015 33544
rect 40957 33535 41015 33541
rect 41322 33532 41328 33544
rect 41380 33572 41386 33584
rect 42613 33575 42671 33581
rect 42613 33572 42625 33575
rect 41380 33544 42625 33572
rect 41380 33532 41386 33544
rect 42613 33541 42625 33544
rect 42659 33541 42671 33575
rect 42613 33535 42671 33541
rect 42705 33575 42763 33581
rect 42705 33541 42717 33575
rect 42751 33572 42763 33575
rect 42812 33572 42840 33600
rect 42751 33544 42840 33572
rect 42751 33541 42763 33544
rect 42705 33535 42763 33541
rect 42886 33532 42892 33584
rect 42944 33572 42950 33584
rect 43901 33575 43959 33581
rect 43901 33572 43913 33575
rect 42944 33544 43913 33572
rect 42944 33532 42950 33544
rect 43901 33541 43913 33544
rect 43947 33541 43959 33575
rect 43901 33535 43959 33541
rect 44117 33575 44175 33581
rect 44117 33541 44129 33575
rect 44163 33572 44175 33575
rect 44358 33572 44364 33584
rect 44163 33544 44364 33572
rect 44163 33541 44175 33544
rect 44117 33535 44175 33541
rect 24118 33504 24124 33516
rect 24079 33476 24124 33504
rect 24118 33464 24124 33476
rect 24176 33464 24182 33516
rect 24765 33507 24823 33513
rect 24765 33473 24777 33507
rect 24811 33504 24823 33507
rect 24854 33504 24860 33516
rect 24811 33476 24860 33504
rect 24811 33473 24823 33476
rect 24765 33467 24823 33473
rect 23937 33439 23995 33445
rect 23937 33405 23949 33439
rect 23983 33436 23995 33439
rect 24026 33436 24032 33448
rect 23983 33408 24032 33436
rect 23983 33405 23995 33408
rect 23937 33399 23995 33405
rect 24026 33396 24032 33408
rect 24084 33436 24090 33448
rect 24780 33436 24808 33467
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 24949 33507 25007 33513
rect 24949 33473 24961 33507
rect 24995 33473 25007 33507
rect 24949 33467 25007 33473
rect 25961 33507 26019 33513
rect 25961 33473 25973 33507
rect 26007 33504 26019 33507
rect 26234 33504 26240 33516
rect 26007 33476 26240 33504
rect 26007 33473 26019 33476
rect 25961 33467 26019 33473
rect 24084 33408 24808 33436
rect 24964 33436 24992 33467
rect 26234 33464 26240 33476
rect 26292 33464 26298 33516
rect 30926 33504 30932 33516
rect 30887 33476 30932 33504
rect 30926 33464 30932 33476
rect 30984 33464 30990 33516
rect 41874 33464 41880 33516
rect 41932 33504 41938 33516
rect 42426 33504 42432 33516
rect 41932 33476 42432 33504
rect 41932 33464 41938 33476
rect 42426 33464 42432 33476
rect 42484 33464 42490 33516
rect 42797 33507 42855 33513
rect 42797 33473 42809 33507
rect 42843 33473 42855 33507
rect 43916 33504 43944 33535
rect 44358 33532 44364 33544
rect 44416 33572 44422 33584
rect 44416 33544 45048 33572
rect 44416 33532 44422 33544
rect 44729 33507 44787 33513
rect 44729 33504 44741 33507
rect 43916 33476 44741 33504
rect 42797 33467 42855 33473
rect 44729 33473 44741 33476
rect 44775 33473 44787 33507
rect 44910 33504 44916 33516
rect 44871 33476 44916 33504
rect 44729 33467 44787 33473
rect 26145 33439 26203 33445
rect 24964 33408 26096 33436
rect 24084 33396 24090 33408
rect 24946 33328 24952 33380
rect 25004 33368 25010 33380
rect 25593 33371 25651 33377
rect 25593 33368 25605 33371
rect 25004 33340 25605 33368
rect 25004 33328 25010 33340
rect 25593 33337 25605 33340
rect 25639 33337 25651 33371
rect 26068 33368 26096 33408
rect 26145 33405 26157 33439
rect 26191 33436 26203 33439
rect 26878 33436 26884 33448
rect 26191 33408 26884 33436
rect 26191 33405 26203 33408
rect 26145 33399 26203 33405
rect 26878 33396 26884 33408
rect 26936 33396 26942 33448
rect 26970 33396 26976 33448
rect 27028 33436 27034 33448
rect 27525 33439 27583 33445
rect 27525 33436 27537 33439
rect 27028 33408 27537 33436
rect 27028 33396 27034 33408
rect 27525 33405 27537 33408
rect 27571 33405 27583 33439
rect 27525 33399 27583 33405
rect 41230 33396 41236 33448
rect 41288 33436 41294 33448
rect 41325 33439 41383 33445
rect 41325 33436 41337 33439
rect 41288 33408 41337 33436
rect 41288 33396 41294 33408
rect 41325 33405 41337 33408
rect 41371 33405 41383 33439
rect 41325 33399 41383 33405
rect 41417 33439 41475 33445
rect 41417 33405 41429 33439
rect 41463 33436 41475 33439
rect 42702 33436 42708 33448
rect 41463 33408 42708 33436
rect 41463 33405 41475 33408
rect 41417 33399 41475 33405
rect 42702 33396 42708 33408
rect 42760 33436 42766 33448
rect 42812 33436 42840 33467
rect 44910 33464 44916 33476
rect 44968 33464 44974 33516
rect 45020 33513 45048 33544
rect 45094 33532 45100 33584
rect 45152 33572 45158 33584
rect 47872 33572 47900 33603
rect 48406 33600 48412 33652
rect 48464 33640 48470 33652
rect 48590 33640 48596 33652
rect 48464 33612 48596 33640
rect 48464 33600 48470 33612
rect 48590 33600 48596 33612
rect 48648 33600 48654 33652
rect 49881 33643 49939 33649
rect 49881 33609 49893 33643
rect 49927 33640 49939 33643
rect 49927 33612 50568 33640
rect 49927 33609 49939 33612
rect 49881 33603 49939 33609
rect 45152 33544 47900 33572
rect 49789 33575 49847 33581
rect 45152 33532 45158 33544
rect 49789 33541 49801 33575
rect 49835 33572 49847 33575
rect 49970 33572 49976 33584
rect 49835 33544 49976 33572
rect 49835 33541 49847 33544
rect 49789 33535 49847 33541
rect 49970 33532 49976 33544
rect 50028 33532 50034 33584
rect 50540 33572 50568 33612
rect 50614 33600 50620 33652
rect 50672 33640 50678 33652
rect 51537 33643 51595 33649
rect 50672 33612 51074 33640
rect 50672 33600 50678 33612
rect 50890 33572 50896 33584
rect 50540 33544 50896 33572
rect 50890 33532 50896 33544
rect 50948 33532 50954 33584
rect 51046 33572 51074 33612
rect 51537 33609 51549 33643
rect 51583 33640 51595 33643
rect 51994 33640 52000 33652
rect 51583 33612 52000 33640
rect 51583 33609 51595 33612
rect 51537 33603 51595 33609
rect 51994 33600 52000 33612
rect 52052 33600 52058 33652
rect 55033 33643 55091 33649
rect 55033 33609 55045 33643
rect 55079 33640 55091 33643
rect 55582 33640 55588 33652
rect 55079 33612 55588 33640
rect 55079 33609 55091 33612
rect 55033 33603 55091 33609
rect 55582 33600 55588 33612
rect 55640 33600 55646 33652
rect 55858 33640 55864 33652
rect 55819 33612 55864 33640
rect 55858 33600 55864 33612
rect 55916 33600 55922 33652
rect 51046 33544 51580 33572
rect 45005 33507 45063 33513
rect 45005 33473 45017 33507
rect 45051 33504 45063 33507
rect 45465 33507 45523 33513
rect 45465 33504 45477 33507
rect 45051 33476 45477 33504
rect 45051 33473 45063 33476
rect 45005 33467 45063 33473
rect 45465 33473 45477 33476
rect 45511 33473 45523 33507
rect 45465 33467 45523 33473
rect 45649 33507 45707 33513
rect 45649 33473 45661 33507
rect 45695 33473 45707 33507
rect 45649 33467 45707 33473
rect 42760 33408 42840 33436
rect 42760 33396 42766 33408
rect 43898 33396 43904 33448
rect 43956 33436 43962 33448
rect 44928 33436 44956 33464
rect 45664 33436 45692 33467
rect 47026 33464 47032 33516
rect 47084 33504 47090 33516
rect 47302 33504 47308 33516
rect 47084 33476 47308 33504
rect 47084 33464 47090 33476
rect 47302 33464 47308 33476
rect 47360 33464 47366 33516
rect 47486 33464 47492 33516
rect 47544 33504 47550 33516
rect 47581 33507 47639 33513
rect 47581 33504 47593 33507
rect 47544 33476 47593 33504
rect 47544 33464 47550 33476
rect 47581 33473 47593 33476
rect 47627 33473 47639 33507
rect 47946 33504 47952 33516
rect 47907 33476 47952 33504
rect 47581 33467 47639 33473
rect 47946 33464 47952 33476
rect 48004 33464 48010 33516
rect 49050 33504 49056 33516
rect 49011 33476 49056 33504
rect 49050 33464 49056 33476
rect 49108 33464 49114 33516
rect 49234 33504 49240 33516
rect 49195 33476 49240 33504
rect 49234 33464 49240 33476
rect 49292 33464 49298 33516
rect 50617 33507 50675 33513
rect 50617 33473 50629 33507
rect 50663 33504 50675 33507
rect 51074 33504 51080 33516
rect 50663 33476 51080 33504
rect 50663 33473 50675 33476
rect 50617 33467 50675 33473
rect 51074 33464 51080 33476
rect 51132 33464 51138 33516
rect 51350 33504 51356 33516
rect 51311 33476 51356 33504
rect 51350 33464 51356 33476
rect 51408 33464 51414 33516
rect 51552 33513 51580 33544
rect 52362 33532 52368 33584
rect 52420 33572 52426 33584
rect 53926 33572 53932 33584
rect 52420 33544 53932 33572
rect 52420 33532 52426 33544
rect 53926 33532 53932 33544
rect 53984 33532 53990 33584
rect 54202 33581 54208 33584
rect 54145 33575 54208 33581
rect 54145 33541 54157 33575
rect 54191 33541 54208 33575
rect 54145 33535 54208 33541
rect 54202 33532 54208 33535
rect 54260 33532 54266 33584
rect 56318 33572 56324 33584
rect 54772 33544 55628 33572
rect 56279 33544 56324 33572
rect 54772 33516 54800 33544
rect 51537 33507 51595 33513
rect 51537 33473 51549 33507
rect 51583 33473 51595 33507
rect 54754 33504 54760 33516
rect 54715 33476 54760 33504
rect 51537 33467 51595 33473
rect 54754 33464 54760 33476
rect 54812 33464 54818 33516
rect 55398 33504 55404 33516
rect 55048 33476 55404 33504
rect 43956 33408 44864 33436
rect 44928 33408 45692 33436
rect 43956 33396 43962 33408
rect 26326 33368 26332 33380
rect 26068 33340 26332 33368
rect 25593 33331 25651 33337
rect 26326 33328 26332 33340
rect 26384 33328 26390 33380
rect 44729 33371 44787 33377
rect 44729 33368 44741 33371
rect 44652 33340 44741 33368
rect 44652 33312 44680 33340
rect 44729 33337 44741 33340
rect 44775 33337 44787 33371
rect 44836 33368 44864 33408
rect 47118 33396 47124 33448
rect 47176 33436 47182 33448
rect 47765 33439 47823 33445
rect 47765 33436 47777 33439
rect 47176 33408 47777 33436
rect 47176 33396 47182 33408
rect 47765 33405 47777 33408
rect 47811 33405 47823 33439
rect 47765 33399 47823 33405
rect 49145 33439 49203 33445
rect 49145 33405 49157 33439
rect 49191 33436 49203 33439
rect 50798 33436 50804 33448
rect 49191 33408 50804 33436
rect 49191 33405 49203 33408
rect 49145 33399 49203 33405
rect 50798 33396 50804 33408
rect 50856 33396 50862 33448
rect 50893 33439 50951 33445
rect 50893 33405 50905 33439
rect 50939 33436 50951 33439
rect 50982 33436 50988 33448
rect 50939 33408 50988 33436
rect 50939 33405 50951 33408
rect 50893 33399 50951 33405
rect 50982 33396 50988 33408
rect 51040 33396 51046 33448
rect 55048 33445 55076 33476
rect 55398 33464 55404 33476
rect 55456 33504 55462 33516
rect 55493 33507 55551 33513
rect 55493 33504 55505 33507
rect 55456 33476 55505 33504
rect 55456 33464 55462 33476
rect 55493 33473 55505 33476
rect 55539 33473 55551 33507
rect 55493 33467 55551 33473
rect 55600 33445 55628 33544
rect 56318 33532 56324 33544
rect 56376 33532 56382 33584
rect 56410 33464 56416 33516
rect 56468 33504 56474 33516
rect 56505 33507 56563 33513
rect 56505 33504 56517 33507
rect 56468 33476 56517 33504
rect 56468 33464 56474 33476
rect 56505 33473 56517 33476
rect 56551 33473 56563 33507
rect 56505 33467 56563 33473
rect 56594 33464 56600 33516
rect 56652 33504 56658 33516
rect 56652 33476 56697 33504
rect 56652 33464 56658 33476
rect 56870 33464 56876 33516
rect 56928 33504 56934 33516
rect 57057 33507 57115 33513
rect 57057 33504 57069 33507
rect 56928 33476 57069 33504
rect 56928 33464 56934 33476
rect 57057 33473 57069 33476
rect 57103 33473 57115 33507
rect 57057 33467 57115 33473
rect 55033 33439 55091 33445
rect 55033 33405 55045 33439
rect 55079 33405 55091 33439
rect 55033 33399 55091 33405
rect 55585 33439 55643 33445
rect 55585 33405 55597 33439
rect 55631 33405 55643 33439
rect 55585 33399 55643 33405
rect 49326 33368 49332 33380
rect 44836 33340 49332 33368
rect 44729 33331 44787 33337
rect 49326 33328 49332 33340
rect 49384 33328 49390 33380
rect 50433 33371 50491 33377
rect 50433 33337 50445 33371
rect 50479 33368 50491 33371
rect 51074 33368 51080 33380
rect 50479 33340 51080 33368
rect 50479 33337 50491 33340
rect 50433 33331 50491 33337
rect 51074 33328 51080 33340
rect 51132 33328 51138 33380
rect 54297 33371 54355 33377
rect 54297 33337 54309 33371
rect 54343 33368 54355 33371
rect 54662 33368 54668 33380
rect 54343 33340 54668 33368
rect 54343 33337 54355 33340
rect 54297 33331 54355 33337
rect 54662 33328 54668 33340
rect 54720 33368 54726 33380
rect 54849 33371 54907 33377
rect 54849 33368 54861 33371
rect 54720 33340 54861 33368
rect 54720 33328 54726 33340
rect 54849 33337 54861 33340
rect 54895 33368 54907 33371
rect 54895 33340 55536 33368
rect 54895 33337 54907 33340
rect 54849 33331 54907 33337
rect 23842 33260 23848 33312
rect 23900 33300 23906 33312
rect 24305 33303 24363 33309
rect 24305 33300 24317 33303
rect 23900 33272 24317 33300
rect 23900 33260 23906 33272
rect 24305 33269 24317 33272
rect 24351 33269 24363 33303
rect 24305 33263 24363 33269
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 27154 33300 27160 33312
rect 25179 33272 27160 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 27154 33260 27160 33272
rect 27212 33260 27218 33312
rect 28905 33303 28963 33309
rect 28905 33269 28917 33303
rect 28951 33300 28963 33303
rect 29086 33300 29092 33312
rect 28951 33272 29092 33300
rect 28951 33269 28963 33272
rect 28905 33263 28963 33269
rect 29086 33260 29092 33272
rect 29144 33260 29150 33312
rect 39114 33260 39120 33312
rect 39172 33300 39178 33312
rect 43898 33300 43904 33312
rect 39172 33272 43904 33300
rect 39172 33260 39178 33272
rect 43898 33260 43904 33272
rect 43956 33260 43962 33312
rect 44085 33303 44143 33309
rect 44085 33269 44097 33303
rect 44131 33300 44143 33303
rect 44174 33300 44180 33312
rect 44131 33272 44180 33300
rect 44131 33269 44143 33272
rect 44085 33263 44143 33269
rect 44174 33260 44180 33272
rect 44232 33260 44238 33312
rect 44634 33260 44640 33312
rect 44692 33260 44698 33312
rect 45554 33260 45560 33312
rect 45612 33300 45618 33312
rect 47578 33300 47584 33312
rect 45612 33272 47584 33300
rect 45612 33260 45618 33272
rect 47578 33260 47584 33272
rect 47636 33260 47642 33312
rect 54110 33300 54116 33312
rect 54071 33272 54116 33300
rect 54110 33260 54116 33272
rect 54168 33260 54174 33312
rect 55508 33309 55536 33340
rect 55493 33303 55551 33309
rect 55493 33269 55505 33303
rect 55539 33269 55551 33303
rect 55493 33263 55551 33269
rect 56321 33303 56379 33309
rect 56321 33269 56333 33303
rect 56367 33300 56379 33303
rect 56962 33300 56968 33312
rect 56367 33272 56968 33300
rect 56367 33269 56379 33272
rect 56321 33263 56379 33269
rect 56962 33260 56968 33272
rect 57020 33260 57026 33312
rect 57146 33300 57152 33312
rect 57107 33272 57152 33300
rect 57146 33260 57152 33272
rect 57204 33260 57210 33312
rect 57238 33260 57244 33312
rect 57296 33300 57302 33312
rect 58069 33303 58127 33309
rect 58069 33300 58081 33303
rect 57296 33272 58081 33300
rect 57296 33260 57302 33272
rect 58069 33269 58081 33272
rect 58115 33269 58127 33303
rect 58069 33263 58127 33269
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 26237 33099 26295 33105
rect 26237 33065 26249 33099
rect 26283 33096 26295 33099
rect 26326 33096 26332 33108
rect 26283 33068 26332 33096
rect 26283 33065 26295 33068
rect 26237 33059 26295 33065
rect 26326 33056 26332 33068
rect 26384 33056 26390 33108
rect 41322 33096 41328 33108
rect 41283 33068 41328 33096
rect 41322 33056 41328 33068
rect 41380 33056 41386 33108
rect 42702 33096 42708 33108
rect 42663 33068 42708 33096
rect 42702 33056 42708 33068
rect 42760 33056 42766 33108
rect 44082 33096 44088 33108
rect 44043 33068 44088 33096
rect 44082 33056 44088 33068
rect 44140 33056 44146 33108
rect 44174 33056 44180 33108
rect 44232 33096 44238 33108
rect 44910 33096 44916 33108
rect 44232 33068 44916 33096
rect 44232 33056 44238 33068
rect 44910 33056 44916 33068
rect 44968 33056 44974 33108
rect 45370 33056 45376 33108
rect 45428 33096 45434 33108
rect 46474 33096 46480 33108
rect 45428 33068 46480 33096
rect 45428 33056 45434 33068
rect 46474 33056 46480 33068
rect 46532 33056 46538 33108
rect 46569 33099 46627 33105
rect 46569 33065 46581 33099
rect 46615 33096 46627 33099
rect 46750 33096 46756 33108
rect 46615 33068 46756 33096
rect 46615 33065 46627 33068
rect 46569 33059 46627 33065
rect 46750 33056 46756 33068
rect 46808 33056 46814 33108
rect 47118 33096 47124 33108
rect 47079 33068 47124 33096
rect 47118 33056 47124 33068
rect 47176 33056 47182 33108
rect 48038 33096 48044 33108
rect 47228 33068 48044 33096
rect 29914 32988 29920 33040
rect 29972 33028 29978 33040
rect 42518 33028 42524 33040
rect 29972 33000 30144 33028
rect 29972 32988 29978 33000
rect 26694 32960 26700 32972
rect 26655 32932 26700 32960
rect 26694 32920 26700 32932
rect 26752 32920 26758 32972
rect 26878 32960 26884 32972
rect 26839 32932 26884 32960
rect 26878 32920 26884 32932
rect 26936 32920 26942 32972
rect 26970 32920 26976 32972
rect 27028 32960 27034 32972
rect 27617 32963 27675 32969
rect 27617 32960 27629 32963
rect 27028 32932 27629 32960
rect 27028 32920 27034 32932
rect 27617 32929 27629 32932
rect 27663 32929 27675 32963
rect 30006 32960 30012 32972
rect 29967 32932 30012 32960
rect 27617 32923 27675 32929
rect 30006 32920 30012 32932
rect 30064 32920 30070 32972
rect 30116 32969 30144 33000
rect 41800 33000 42524 33028
rect 30101 32963 30159 32969
rect 30101 32929 30113 32963
rect 30147 32960 30159 32963
rect 30282 32960 30288 32972
rect 30147 32932 30288 32960
rect 30147 32929 30159 32932
rect 30101 32923 30159 32929
rect 30282 32920 30288 32932
rect 30340 32920 30346 32972
rect 23842 32892 23848 32904
rect 23803 32864 23848 32892
rect 23842 32852 23848 32864
rect 23900 32852 23906 32904
rect 24397 32895 24455 32901
rect 24397 32861 24409 32895
rect 24443 32892 24455 32895
rect 25038 32892 25044 32904
rect 24443 32864 25044 32892
rect 24443 32861 24455 32864
rect 24397 32855 24455 32861
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 35802 32852 35808 32904
rect 35860 32892 35866 32904
rect 37090 32901 37096 32904
rect 36817 32895 36875 32901
rect 36817 32892 36829 32895
rect 35860 32864 36829 32892
rect 35860 32852 35866 32864
rect 36817 32861 36829 32864
rect 36863 32861 36875 32895
rect 37084 32892 37096 32901
rect 37051 32864 37096 32892
rect 36817 32855 36875 32861
rect 37084 32855 37096 32864
rect 37090 32852 37096 32855
rect 37148 32852 37154 32904
rect 41506 32892 41512 32904
rect 41467 32864 41512 32892
rect 41506 32852 41512 32864
rect 41564 32852 41570 32904
rect 41598 32852 41604 32904
rect 41656 32892 41662 32904
rect 41800 32901 41828 33000
rect 42518 32988 42524 33000
rect 42576 33028 42582 33040
rect 47228 33028 47256 33068
rect 48038 33056 48044 33068
rect 48096 33056 48102 33108
rect 48130 33056 48136 33108
rect 48188 33096 48194 33108
rect 48225 33099 48283 33105
rect 48225 33096 48237 33099
rect 48188 33068 48237 33096
rect 48188 33056 48194 33068
rect 48225 33065 48237 33068
rect 48271 33065 48283 33099
rect 48225 33059 48283 33065
rect 50154 33056 50160 33108
rect 50212 33096 50218 33108
rect 51077 33099 51135 33105
rect 51077 33096 51089 33099
rect 50212 33068 51089 33096
rect 50212 33056 50218 33068
rect 51077 33065 51089 33068
rect 51123 33096 51135 33099
rect 51350 33096 51356 33108
rect 51123 33068 51356 33096
rect 51123 33065 51135 33068
rect 51077 33059 51135 33065
rect 51350 33056 51356 33068
rect 51408 33056 51414 33108
rect 53837 33099 53895 33105
rect 53837 33065 53849 33099
rect 53883 33096 53895 33099
rect 54478 33096 54484 33108
rect 53883 33068 54484 33096
rect 53883 33065 53895 33068
rect 53837 33059 53895 33065
rect 54478 33056 54484 33068
rect 54536 33056 54542 33108
rect 55582 33056 55588 33108
rect 55640 33096 55646 33108
rect 55677 33099 55735 33105
rect 55677 33096 55689 33099
rect 55640 33068 55689 33096
rect 55640 33056 55646 33068
rect 55677 33065 55689 33068
rect 55723 33096 55735 33099
rect 56410 33096 56416 33108
rect 55723 33068 56416 33096
rect 55723 33065 55735 33068
rect 55677 33059 55735 33065
rect 56410 33056 56416 33068
rect 56468 33056 56474 33108
rect 42576 33000 47256 33028
rect 42576 32988 42582 33000
rect 44450 32960 44456 32972
rect 44100 32932 44456 32960
rect 44100 32901 44128 32932
rect 44450 32920 44456 32932
rect 44508 32920 44514 32972
rect 41785 32895 41843 32901
rect 41656 32864 41701 32892
rect 41656 32852 41662 32864
rect 41785 32861 41797 32895
rect 41831 32861 41843 32895
rect 41785 32855 41843 32861
rect 41877 32895 41935 32901
rect 41877 32861 41889 32895
rect 41923 32892 41935 32895
rect 44085 32895 44143 32901
rect 41923 32864 42564 32892
rect 41923 32861 41935 32864
rect 41877 32855 41935 32861
rect 24642 32827 24700 32833
rect 24642 32824 24654 32827
rect 23676 32796 24654 32824
rect 23676 32765 23704 32796
rect 24642 32793 24654 32796
rect 24688 32793 24700 32827
rect 24642 32787 24700 32793
rect 27884 32827 27942 32833
rect 27884 32793 27896 32827
rect 27930 32824 27942 32827
rect 28534 32824 28540 32836
rect 27930 32796 28540 32824
rect 27930 32793 27942 32796
rect 27884 32787 27942 32793
rect 28534 32784 28540 32796
rect 28592 32784 28598 32836
rect 29917 32827 29975 32833
rect 29917 32824 29929 32827
rect 29012 32796 29929 32824
rect 29012 32768 29040 32796
rect 29917 32793 29929 32796
rect 29963 32793 29975 32827
rect 29917 32787 29975 32793
rect 41230 32784 41236 32836
rect 41288 32824 41294 32836
rect 41892 32824 41920 32855
rect 42536 32833 42564 32864
rect 44085 32861 44097 32895
rect 44131 32861 44143 32895
rect 44085 32855 44143 32861
rect 44269 32895 44327 32901
rect 44269 32861 44281 32895
rect 44315 32892 44327 32895
rect 44818 32892 44824 32904
rect 44315 32864 44824 32892
rect 44315 32861 44327 32864
rect 44269 32855 44327 32861
rect 44818 32852 44824 32864
rect 44876 32852 44882 32904
rect 45278 32852 45284 32904
rect 45336 32892 45342 32904
rect 45664 32901 45692 33000
rect 47946 32988 47952 33040
rect 48004 33028 48010 33040
rect 48409 33031 48467 33037
rect 48409 33028 48421 33031
rect 48004 33000 48421 33028
rect 48004 32988 48010 33000
rect 48409 32997 48421 33000
rect 48455 32997 48467 33031
rect 51258 33028 51264 33040
rect 51219 33000 51264 33028
rect 48409 32991 48467 32997
rect 51258 32988 51264 33000
rect 51316 32988 51322 33040
rect 46492 32932 47716 32960
rect 45465 32895 45523 32901
rect 45465 32892 45477 32895
rect 45336 32864 45477 32892
rect 45336 32852 45342 32864
rect 45465 32861 45477 32864
rect 45511 32861 45523 32895
rect 45465 32855 45523 32861
rect 45649 32895 45707 32901
rect 45649 32861 45661 32895
rect 45695 32861 45707 32895
rect 45649 32855 45707 32861
rect 46382 32852 46388 32904
rect 46440 32892 46446 32904
rect 46492 32901 46520 32932
rect 46477 32895 46535 32901
rect 46477 32892 46489 32895
rect 46440 32864 46489 32892
rect 46440 32852 46446 32864
rect 46477 32861 46489 32864
rect 46523 32861 46535 32895
rect 46477 32855 46535 32861
rect 46661 32895 46719 32901
rect 46661 32861 46673 32895
rect 46707 32892 46719 32895
rect 47305 32895 47363 32901
rect 46707 32864 47256 32892
rect 46707 32861 46719 32864
rect 46661 32855 46719 32861
rect 41288 32796 41920 32824
rect 42337 32827 42395 32833
rect 41288 32784 41294 32796
rect 42337 32793 42349 32827
rect 42383 32793 42395 32827
rect 42337 32787 42395 32793
rect 42521 32827 42579 32833
rect 42521 32793 42533 32827
rect 42567 32824 42579 32827
rect 42567 32796 44312 32824
rect 42567 32793 42579 32796
rect 42521 32787 42579 32793
rect 23661 32759 23719 32765
rect 23661 32725 23673 32759
rect 23707 32725 23719 32759
rect 23661 32719 23719 32725
rect 25777 32759 25835 32765
rect 25777 32725 25789 32759
rect 25823 32756 25835 32759
rect 26050 32756 26056 32768
rect 25823 32728 26056 32756
rect 25823 32725 25835 32728
rect 25777 32719 25835 32725
rect 26050 32716 26056 32728
rect 26108 32716 26114 32768
rect 26605 32759 26663 32765
rect 26605 32725 26617 32759
rect 26651 32756 26663 32759
rect 27982 32756 27988 32768
rect 26651 32728 27988 32756
rect 26651 32725 26663 32728
rect 26605 32719 26663 32725
rect 27982 32716 27988 32728
rect 28040 32716 28046 32768
rect 28994 32756 29000 32768
rect 28955 32728 29000 32756
rect 28994 32716 29000 32728
rect 29052 32716 29058 32768
rect 29546 32756 29552 32768
rect 29507 32728 29552 32756
rect 29546 32716 29552 32728
rect 29604 32716 29610 32768
rect 38197 32759 38255 32765
rect 38197 32725 38209 32759
rect 38243 32756 38255 32759
rect 38746 32756 38752 32768
rect 38243 32728 38752 32756
rect 38243 32725 38255 32728
rect 38197 32719 38255 32725
rect 38746 32716 38752 32728
rect 38804 32716 38810 32768
rect 41598 32716 41604 32768
rect 41656 32756 41662 32768
rect 42352 32756 42380 32787
rect 44284 32768 44312 32796
rect 42610 32756 42616 32768
rect 41656 32728 42616 32756
rect 41656 32716 41662 32728
rect 42610 32716 42616 32728
rect 42668 32716 42674 32768
rect 44266 32716 44272 32768
rect 44324 32716 44330 32768
rect 45186 32716 45192 32768
rect 45244 32756 45250 32768
rect 45557 32759 45615 32765
rect 45557 32756 45569 32759
rect 45244 32728 45569 32756
rect 45244 32716 45250 32728
rect 45557 32725 45569 32728
rect 45603 32725 45615 32759
rect 47228 32756 47256 32864
rect 47305 32861 47317 32895
rect 47351 32892 47363 32895
rect 47486 32892 47492 32904
rect 47351 32864 47492 32892
rect 47351 32861 47363 32864
rect 47305 32855 47363 32861
rect 47486 32852 47492 32864
rect 47544 32852 47550 32904
rect 47581 32895 47639 32901
rect 47581 32861 47593 32895
rect 47627 32892 47639 32895
rect 47688 32892 47716 32932
rect 47854 32920 47860 32972
rect 47912 32960 47918 32972
rect 50062 32960 50068 32972
rect 47912 32932 50068 32960
rect 47912 32920 47918 32932
rect 50062 32920 50068 32932
rect 50120 32960 50126 32972
rect 50433 32963 50491 32969
rect 50433 32960 50445 32963
rect 50120 32932 50445 32960
rect 50120 32920 50126 32932
rect 50433 32929 50445 32932
rect 50479 32929 50491 32963
rect 51368 32960 51396 33056
rect 51721 33031 51779 33037
rect 51721 32997 51733 33031
rect 51767 33028 51779 33031
rect 51810 33028 51816 33040
rect 51767 33000 51816 33028
rect 51767 32997 51779 33000
rect 51721 32991 51779 32997
rect 51810 32988 51816 33000
rect 51868 32988 51874 33040
rect 57238 33028 57244 33040
rect 56336 33000 57244 33028
rect 56336 32969 56364 33000
rect 57238 32988 57244 33000
rect 57296 32988 57302 33040
rect 56321 32963 56379 32969
rect 51368 32932 52040 32960
rect 50433 32923 50491 32929
rect 47627 32867 48314 32892
rect 47627 32864 48329 32867
rect 47627 32861 47639 32864
rect 47581 32855 47639 32861
rect 48271 32861 48329 32864
rect 47504 32824 47532 32852
rect 48041 32827 48099 32833
rect 48041 32824 48053 32827
rect 47504 32796 48053 32824
rect 48041 32793 48053 32796
rect 48087 32793 48099 32827
rect 48271 32827 48283 32861
rect 48317 32827 48329 32861
rect 48271 32821 48329 32827
rect 48041 32787 48099 32793
rect 47489 32759 47547 32765
rect 47489 32756 47501 32759
rect 47228 32728 47501 32756
rect 45557 32719 45615 32725
rect 47489 32725 47501 32728
rect 47535 32756 47547 32759
rect 47946 32756 47952 32768
rect 47535 32728 47952 32756
rect 47535 32725 47547 32728
rect 47489 32719 47547 32725
rect 47946 32716 47952 32728
rect 48004 32716 48010 32768
rect 48056 32756 48084 32787
rect 49234 32784 49240 32836
rect 49292 32824 49298 32836
rect 50154 32824 50160 32836
rect 49292 32796 50160 32824
rect 49292 32784 49298 32796
rect 50154 32784 50160 32796
rect 50212 32824 50218 32836
rect 50249 32827 50307 32833
rect 50249 32824 50261 32827
rect 50212 32796 50261 32824
rect 50212 32784 50218 32796
rect 50249 32793 50261 32796
rect 50295 32793 50307 32827
rect 50249 32787 50307 32793
rect 49602 32756 49608 32768
rect 48056 32728 49608 32756
rect 49602 32716 49608 32728
rect 49660 32716 49666 32768
rect 50448 32756 50476 32923
rect 52012 32901 52040 32932
rect 56321 32929 56333 32963
rect 56367 32929 56379 32963
rect 56321 32923 56379 32929
rect 56505 32963 56563 32969
rect 56505 32929 56517 32963
rect 56551 32960 56563 32963
rect 57146 32960 57152 32972
rect 56551 32932 57152 32960
rect 56551 32929 56563 32932
rect 56505 32923 56563 32929
rect 57146 32920 57152 32932
rect 57204 32920 57210 32972
rect 57790 32960 57796 32972
rect 57751 32932 57796 32960
rect 57790 32920 57796 32932
rect 57848 32920 57854 32972
rect 51905 32895 51963 32901
rect 51905 32892 51917 32895
rect 50908 32864 51917 32892
rect 50908 32836 50936 32864
rect 51905 32861 51917 32864
rect 51951 32861 51963 32895
rect 51905 32855 51963 32861
rect 51997 32895 52055 32901
rect 51997 32861 52009 32895
rect 52043 32861 52055 32895
rect 54110 32892 54116 32904
rect 51997 32855 52055 32861
rect 53116 32864 54116 32892
rect 50890 32824 50896 32836
rect 50851 32796 50896 32824
rect 50890 32784 50896 32796
rect 50948 32784 50954 32836
rect 51074 32784 51080 32836
rect 51132 32833 51138 32836
rect 51132 32827 51151 32833
rect 51139 32824 51151 32827
rect 51721 32827 51779 32833
rect 51721 32824 51733 32827
rect 51139 32796 51733 32824
rect 51139 32793 51151 32796
rect 51132 32787 51151 32793
rect 51721 32793 51733 32796
rect 51767 32793 51779 32827
rect 51721 32787 51779 32793
rect 51132 32784 51138 32787
rect 53116 32756 53144 32864
rect 54110 32852 54116 32864
rect 54168 32852 54174 32904
rect 54570 32892 54576 32904
rect 54531 32864 54576 32892
rect 54570 32852 54576 32864
rect 54628 32852 54634 32904
rect 54754 32892 54760 32904
rect 54715 32864 54760 32892
rect 54754 32852 54760 32864
rect 54812 32852 54818 32904
rect 53837 32827 53895 32833
rect 53837 32793 53849 32827
rect 53883 32824 53895 32827
rect 54202 32824 54208 32836
rect 53883 32796 54208 32824
rect 53883 32793 53895 32796
rect 53837 32787 53895 32793
rect 54202 32784 54208 32796
rect 54260 32824 54266 32836
rect 54665 32827 54723 32833
rect 54665 32824 54677 32827
rect 54260 32796 54677 32824
rect 54260 32784 54266 32796
rect 54665 32793 54677 32796
rect 54711 32793 54723 32827
rect 55490 32824 55496 32836
rect 55451 32796 55496 32824
rect 54665 32787 54723 32793
rect 55490 32784 55496 32796
rect 55548 32784 55554 32836
rect 55709 32827 55767 32833
rect 55709 32793 55721 32827
rect 55755 32824 55767 32827
rect 56594 32824 56600 32836
rect 55755 32796 56600 32824
rect 55755 32793 55767 32796
rect 55709 32787 55767 32793
rect 56594 32784 56600 32796
rect 56652 32784 56658 32836
rect 50448 32728 53144 32756
rect 53926 32716 53932 32768
rect 53984 32756 53990 32768
rect 54021 32759 54079 32765
rect 54021 32756 54033 32759
rect 53984 32728 54033 32756
rect 53984 32716 53990 32728
rect 54021 32725 54033 32728
rect 54067 32725 54079 32759
rect 54021 32719 54079 32725
rect 55861 32759 55919 32765
rect 55861 32725 55873 32759
rect 55907 32756 55919 32759
rect 57146 32756 57152 32768
rect 55907 32728 57152 32756
rect 55907 32725 55919 32728
rect 55861 32719 55919 32725
rect 57146 32716 57152 32728
rect 57204 32716 57210 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 25038 32512 25044 32564
rect 25096 32512 25102 32564
rect 26234 32552 26240 32564
rect 26195 32524 26240 32552
rect 26234 32512 26240 32524
rect 26292 32512 26298 32564
rect 40678 32512 40684 32564
rect 40736 32552 40742 32564
rect 41049 32555 41107 32561
rect 41049 32552 41061 32555
rect 40736 32524 41061 32552
rect 40736 32512 40742 32524
rect 41049 32521 41061 32524
rect 41095 32521 41107 32555
rect 41049 32515 41107 32521
rect 41417 32555 41475 32561
rect 41417 32521 41429 32555
rect 41463 32552 41475 32555
rect 41598 32552 41604 32564
rect 41463 32524 41604 32552
rect 41463 32521 41475 32524
rect 41417 32515 41475 32521
rect 41598 32512 41604 32524
rect 41656 32512 41662 32564
rect 42426 32552 42432 32564
rect 42387 32524 42432 32552
rect 42426 32512 42432 32524
rect 42484 32512 42490 32564
rect 47394 32512 47400 32564
rect 47452 32552 47458 32564
rect 47673 32555 47731 32561
rect 47673 32552 47685 32555
rect 47452 32524 47685 32552
rect 47452 32512 47458 32524
rect 47673 32521 47685 32524
rect 47719 32521 47731 32555
rect 48314 32552 48320 32564
rect 47673 32515 47731 32521
rect 47780 32524 48320 32552
rect 24946 32484 24952 32496
rect 24228 32456 24952 32484
rect 24026 32416 24032 32428
rect 23987 32388 24032 32416
rect 24026 32376 24032 32388
rect 24084 32376 24090 32428
rect 24228 32425 24256 32456
rect 24946 32444 24952 32456
rect 25004 32444 25010 32496
rect 24213 32419 24271 32425
rect 24213 32385 24225 32419
rect 24259 32385 24271 32419
rect 24213 32379 24271 32385
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32416 24915 32419
rect 25056 32416 25084 32512
rect 34698 32484 34704 32496
rect 34164 32456 34704 32484
rect 25130 32425 25136 32428
rect 24903 32388 25084 32416
rect 24903 32385 24915 32388
rect 24857 32379 24915 32385
rect 25124 32379 25136 32425
rect 25188 32416 25194 32428
rect 27154 32416 27160 32428
rect 25188 32388 25224 32416
rect 27115 32388 27160 32416
rect 25130 32376 25136 32379
rect 25188 32376 25194 32388
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 28813 32419 28871 32425
rect 28813 32385 28825 32419
rect 28859 32416 28871 32419
rect 29546 32416 29552 32428
rect 28859 32388 29552 32416
rect 28859 32385 28871 32388
rect 28813 32379 28871 32385
rect 29546 32376 29552 32388
rect 29604 32376 29610 32428
rect 32306 32416 32312 32428
rect 32267 32388 32312 32416
rect 32306 32376 32312 32388
rect 32364 32376 32370 32428
rect 34164 32425 34192 32456
rect 34698 32444 34704 32456
rect 34756 32444 34762 32496
rect 36722 32444 36728 32496
rect 36780 32484 36786 32496
rect 37522 32487 37580 32493
rect 37522 32484 37534 32487
rect 36780 32456 37534 32484
rect 36780 32444 36786 32456
rect 37522 32453 37534 32456
rect 37568 32453 37580 32487
rect 37522 32447 37580 32453
rect 41690 32444 41696 32496
rect 41748 32484 41754 32496
rect 47780 32484 47808 32524
rect 48314 32512 48320 32524
rect 48372 32512 48378 32564
rect 52733 32555 52791 32561
rect 48700 32524 51120 32552
rect 48700 32496 48728 32524
rect 48682 32484 48688 32496
rect 41748 32456 47808 32484
rect 47872 32456 48452 32484
rect 48595 32456 48688 32484
rect 41748 32444 41754 32456
rect 34149 32419 34207 32425
rect 34149 32385 34161 32419
rect 34195 32385 34207 32419
rect 34149 32379 34207 32385
rect 34416 32419 34474 32425
rect 34416 32385 34428 32419
rect 34462 32416 34474 32419
rect 34790 32416 34796 32428
rect 34462 32388 34796 32416
rect 34462 32385 34474 32388
rect 34416 32379 34474 32385
rect 34790 32376 34796 32388
rect 34848 32376 34854 32428
rect 35710 32376 35716 32428
rect 35768 32416 35774 32428
rect 37182 32416 37188 32428
rect 35768 32388 37188 32416
rect 35768 32376 35774 32388
rect 37182 32376 37188 32388
rect 37240 32416 37246 32428
rect 37277 32419 37335 32425
rect 37277 32416 37289 32419
rect 37240 32388 37289 32416
rect 37240 32376 37246 32388
rect 37277 32385 37289 32388
rect 37323 32385 37335 32419
rect 41230 32416 41236 32428
rect 41191 32388 41236 32416
rect 37277 32379 37335 32385
rect 41230 32376 41236 32388
rect 41288 32376 41294 32428
rect 41506 32376 41512 32428
rect 41564 32416 41570 32428
rect 41874 32416 41880 32428
rect 41564 32388 41880 32416
rect 41564 32376 41570 32388
rect 41874 32376 41880 32388
rect 41932 32376 41938 32428
rect 42242 32376 42248 32428
rect 42300 32416 42306 32428
rect 42613 32419 42671 32425
rect 42613 32416 42625 32419
rect 42300 32388 42625 32416
rect 42300 32376 42306 32388
rect 42613 32385 42625 32388
rect 42659 32385 42671 32419
rect 42613 32379 42671 32385
rect 42702 32376 42708 32428
rect 42760 32416 42766 32428
rect 42889 32419 42947 32425
rect 42760 32388 42805 32416
rect 42760 32376 42766 32388
rect 42889 32385 42901 32419
rect 42935 32385 42947 32419
rect 42889 32379 42947 32385
rect 42981 32419 43039 32425
rect 42981 32385 42993 32419
rect 43027 32416 43039 32419
rect 44450 32416 44456 32428
rect 43027 32388 44456 32416
rect 43027 32385 43039 32388
rect 42981 32379 43039 32385
rect 27614 32308 27620 32360
rect 27672 32348 27678 32360
rect 28629 32351 28687 32357
rect 28629 32348 28641 32351
rect 27672 32320 28641 32348
rect 27672 32308 27678 32320
rect 28629 32317 28641 32320
rect 28675 32348 28687 32351
rect 30374 32348 30380 32360
rect 28675 32320 30380 32348
rect 28675 32317 28687 32320
rect 28629 32311 28687 32317
rect 30374 32308 30380 32320
rect 30432 32348 30438 32360
rect 32125 32351 32183 32357
rect 32125 32348 32137 32351
rect 30432 32320 32137 32348
rect 30432 32308 30438 32320
rect 32125 32317 32137 32320
rect 32171 32317 32183 32351
rect 42904 32348 42932 32379
rect 44450 32376 44456 32388
rect 44508 32376 44514 32428
rect 45002 32416 45008 32428
rect 44963 32388 45008 32416
rect 45002 32376 45008 32388
rect 45060 32376 45066 32428
rect 45186 32416 45192 32428
rect 45147 32388 45192 32416
rect 45186 32376 45192 32388
rect 45244 32376 45250 32428
rect 47872 32425 47900 32456
rect 47857 32419 47915 32425
rect 47857 32385 47869 32419
rect 47903 32385 47915 32419
rect 47857 32379 47915 32385
rect 47949 32419 48007 32425
rect 47949 32385 47961 32419
rect 47995 32385 48007 32419
rect 47949 32379 48007 32385
rect 43070 32348 43076 32360
rect 42904 32320 43076 32348
rect 32125 32311 32183 32317
rect 43070 32308 43076 32320
rect 43128 32308 43134 32360
rect 47964 32348 47992 32379
rect 48038 32376 48044 32428
rect 48096 32416 48102 32428
rect 48133 32419 48191 32425
rect 48133 32416 48145 32419
rect 48096 32388 48145 32416
rect 48096 32376 48102 32388
rect 48133 32385 48145 32388
rect 48179 32385 48191 32419
rect 48133 32379 48191 32385
rect 48222 32376 48228 32428
rect 48280 32416 48286 32428
rect 48280 32388 48325 32416
rect 48280 32376 48286 32388
rect 48424 32348 48452 32456
rect 48682 32444 48688 32456
rect 48740 32444 48746 32496
rect 51092 32493 51120 32524
rect 52733 32521 52745 32555
rect 52779 32521 52791 32555
rect 52733 32515 52791 32521
rect 53561 32555 53619 32561
rect 53561 32521 53573 32555
rect 53607 32552 53619 32555
rect 53742 32552 53748 32564
rect 53607 32524 53748 32552
rect 53607 32521 53619 32524
rect 53561 32515 53619 32521
rect 51077 32487 51135 32493
rect 51077 32453 51089 32487
rect 51123 32484 51135 32487
rect 51534 32484 51540 32496
rect 51123 32456 51540 32484
rect 51123 32453 51135 32456
rect 51077 32447 51135 32453
rect 51534 32444 51540 32456
rect 51592 32444 51598 32496
rect 51810 32484 51816 32496
rect 51771 32456 51816 32484
rect 51810 32444 51816 32456
rect 51868 32444 51874 32496
rect 52748 32484 52776 32515
rect 53742 32512 53748 32524
rect 53800 32512 53806 32564
rect 56502 32552 56508 32564
rect 56463 32524 56508 32552
rect 56502 32512 56508 32524
rect 56560 32512 56566 32564
rect 57054 32552 57060 32564
rect 57015 32524 57060 32552
rect 57054 32512 57060 32524
rect 57112 32512 57118 32564
rect 52748 32456 53512 32484
rect 48866 32416 48872 32428
rect 48827 32388 48872 32416
rect 48866 32376 48872 32388
rect 48924 32376 48930 32428
rect 49973 32419 50031 32425
rect 49973 32385 49985 32419
rect 50019 32385 50031 32419
rect 49973 32379 50031 32385
rect 49053 32351 49111 32357
rect 49053 32348 49065 32351
rect 47964 32320 48084 32348
rect 48424 32320 49065 32348
rect 44450 32240 44456 32292
rect 44508 32280 44514 32292
rect 47854 32280 47860 32292
rect 44508 32252 47860 32280
rect 44508 32240 44514 32252
rect 47854 32240 47860 32252
rect 47912 32240 47918 32292
rect 24397 32215 24455 32221
rect 24397 32181 24409 32215
rect 24443 32212 24455 32215
rect 25222 32212 25228 32224
rect 24443 32184 25228 32212
rect 24443 32181 24455 32184
rect 24397 32175 24455 32181
rect 25222 32172 25228 32184
rect 25280 32172 25286 32224
rect 25498 32172 25504 32224
rect 25556 32212 25562 32224
rect 26973 32215 27031 32221
rect 26973 32212 26985 32215
rect 25556 32184 26985 32212
rect 25556 32172 25562 32184
rect 26973 32181 26985 32184
rect 27019 32181 27031 32215
rect 26973 32175 27031 32181
rect 28718 32172 28724 32224
rect 28776 32212 28782 32224
rect 28997 32215 29055 32221
rect 28997 32212 29009 32215
rect 28776 32184 29009 32212
rect 28776 32172 28782 32184
rect 28997 32181 29009 32184
rect 29043 32181 29055 32215
rect 28997 32175 29055 32181
rect 31754 32172 31760 32224
rect 31812 32212 31818 32224
rect 32493 32215 32551 32221
rect 32493 32212 32505 32215
rect 31812 32184 32505 32212
rect 31812 32172 31818 32184
rect 32493 32181 32505 32184
rect 32539 32181 32551 32215
rect 32493 32175 32551 32181
rect 35529 32215 35587 32221
rect 35529 32181 35541 32215
rect 35575 32212 35587 32215
rect 36722 32212 36728 32224
rect 35575 32184 36728 32212
rect 35575 32181 35587 32184
rect 35529 32175 35587 32181
rect 36722 32172 36728 32184
rect 36780 32172 36786 32224
rect 38654 32212 38660 32224
rect 38615 32184 38660 32212
rect 38654 32172 38660 32184
rect 38712 32172 38718 32224
rect 44818 32172 44824 32224
rect 44876 32212 44882 32224
rect 45097 32215 45155 32221
rect 45097 32212 45109 32215
rect 44876 32184 45109 32212
rect 44876 32172 44882 32184
rect 45097 32181 45109 32184
rect 45143 32181 45155 32215
rect 48056 32212 48084 32320
rect 49053 32317 49065 32320
rect 49099 32317 49111 32351
rect 49988 32348 50016 32379
rect 50062 32376 50068 32428
rect 50120 32416 50126 32428
rect 50157 32419 50215 32425
rect 50157 32416 50169 32419
rect 50120 32388 50169 32416
rect 50120 32376 50126 32388
rect 50157 32385 50169 32388
rect 50203 32385 50215 32419
rect 50890 32416 50896 32428
rect 50851 32388 50896 32416
rect 50157 32379 50215 32385
rect 50890 32376 50896 32388
rect 50948 32376 50954 32428
rect 51258 32376 51264 32428
rect 51316 32416 51322 32428
rect 51997 32419 52055 32425
rect 51997 32416 52009 32419
rect 51316 32388 52009 32416
rect 51316 32376 51322 32388
rect 51997 32385 52009 32388
rect 52043 32385 52055 32419
rect 51997 32379 52055 32385
rect 52638 32376 52644 32428
rect 52696 32416 52702 32428
rect 53484 32425 53512 32456
rect 52733 32419 52791 32425
rect 52733 32416 52745 32419
rect 52696 32388 52745 32416
rect 52696 32376 52702 32388
rect 52733 32385 52745 32388
rect 52779 32385 52791 32419
rect 52733 32379 52791 32385
rect 53469 32419 53527 32425
rect 53469 32385 53481 32419
rect 53515 32416 53527 32419
rect 53558 32416 53564 32428
rect 53515 32388 53564 32416
rect 53515 32385 53527 32388
rect 53469 32379 53527 32385
rect 53558 32376 53564 32388
rect 53616 32376 53622 32428
rect 53653 32419 53711 32425
rect 53653 32385 53665 32419
rect 53699 32385 53711 32419
rect 53653 32379 53711 32385
rect 50908 32348 50936 32376
rect 49988 32320 50936 32348
rect 49053 32311 49111 32317
rect 52546 32308 52552 32360
rect 52604 32348 52610 32360
rect 53009 32351 53067 32357
rect 53009 32348 53021 32351
rect 52604 32320 53021 32348
rect 52604 32308 52610 32320
rect 53009 32317 53021 32320
rect 53055 32317 53067 32351
rect 53009 32311 53067 32317
rect 53098 32308 53104 32360
rect 53156 32348 53162 32360
rect 53668 32348 53696 32379
rect 55490 32376 55496 32428
rect 55548 32416 55554 32428
rect 56229 32419 56287 32425
rect 56229 32416 56241 32419
rect 55548 32388 56241 32416
rect 55548 32376 55554 32388
rect 56229 32385 56241 32388
rect 56275 32385 56287 32419
rect 56962 32416 56968 32428
rect 56923 32388 56968 32416
rect 56229 32379 56287 32385
rect 56962 32376 56968 32388
rect 57020 32376 57026 32428
rect 57146 32416 57152 32428
rect 57107 32388 57152 32416
rect 57146 32376 57152 32388
rect 57204 32376 57210 32428
rect 53156 32320 53696 32348
rect 53156 32308 53162 32320
rect 55582 32308 55588 32360
rect 55640 32348 55646 32360
rect 55861 32351 55919 32357
rect 55861 32348 55873 32351
rect 55640 32320 55873 32348
rect 55640 32308 55646 32320
rect 55861 32317 55873 32320
rect 55907 32317 55919 32351
rect 55861 32311 55919 32317
rect 56321 32351 56379 32357
rect 56321 32317 56333 32351
rect 56367 32348 56379 32351
rect 56594 32348 56600 32360
rect 56367 32320 56600 32348
rect 56367 32317 56379 32320
rect 56321 32311 56379 32317
rect 56594 32308 56600 32320
rect 56652 32308 56658 32360
rect 49970 32280 49976 32292
rect 48286 32252 49976 32280
rect 48286 32212 48314 32252
rect 49970 32240 49976 32252
rect 50028 32280 50034 32292
rect 50065 32283 50123 32289
rect 50065 32280 50077 32283
rect 50028 32252 50077 32280
rect 50028 32240 50034 32252
rect 50065 32249 50077 32252
rect 50111 32249 50123 32283
rect 52822 32280 52828 32292
rect 52783 32252 52828 32280
rect 50065 32243 50123 32249
rect 52822 32240 52828 32252
rect 52880 32240 52886 32292
rect 54662 32280 54668 32292
rect 53392 32252 54668 32280
rect 48056 32184 48314 32212
rect 52181 32215 52239 32221
rect 45097 32175 45155 32181
rect 52181 32181 52193 32215
rect 52227 32212 52239 32215
rect 53392 32212 53420 32252
rect 54662 32240 54668 32252
rect 54720 32240 54726 32292
rect 52227 32184 53420 32212
rect 52227 32181 52239 32184
rect 52181 32175 52239 32181
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 28534 32008 28540 32020
rect 28495 31980 28540 32008
rect 28534 31968 28540 31980
rect 28592 31968 28598 32020
rect 32953 32011 33011 32017
rect 32953 32008 32965 32011
rect 31128 31980 32965 32008
rect 26421 31943 26479 31949
rect 26421 31909 26433 31943
rect 26467 31940 26479 31943
rect 27982 31940 27988 31952
rect 26467 31912 27988 31940
rect 26467 31909 26479 31912
rect 26421 31903 26479 31909
rect 27982 31900 27988 31912
rect 28040 31900 28046 31952
rect 25038 31872 25044 31884
rect 24999 31844 25044 31872
rect 25038 31832 25044 31844
rect 25096 31832 25102 31884
rect 30285 31875 30343 31881
rect 30285 31841 30297 31875
rect 30331 31872 30343 31875
rect 30374 31872 30380 31884
rect 30331 31844 30380 31872
rect 30331 31841 30343 31844
rect 30285 31835 30343 31841
rect 30374 31832 30380 31844
rect 30432 31832 30438 31884
rect 30926 31872 30932 31884
rect 30484 31844 30932 31872
rect 25056 31804 25084 31832
rect 26970 31804 26976 31816
rect 25056 31776 26976 31804
rect 26970 31764 26976 31776
rect 27028 31764 27034 31816
rect 28718 31804 28724 31816
rect 28679 31776 28724 31804
rect 28718 31764 28724 31776
rect 28776 31764 28782 31816
rect 30484 31813 30512 31844
rect 30926 31832 30932 31844
rect 30984 31832 30990 31884
rect 31128 31872 31156 31980
rect 32953 31977 32965 31980
rect 32999 31977 33011 32011
rect 32953 31971 33011 31977
rect 41414 31968 41420 32020
rect 41472 32008 41478 32020
rect 41785 32011 41843 32017
rect 41785 32008 41797 32011
rect 41472 31980 41797 32008
rect 41472 31968 41478 31980
rect 41785 31977 41797 31980
rect 41831 31977 41843 32011
rect 41785 31971 41843 31977
rect 42702 31968 42708 32020
rect 42760 32008 42766 32020
rect 42889 32011 42947 32017
rect 42889 32008 42901 32011
rect 42760 31980 42901 32008
rect 42760 31968 42766 31980
rect 42889 31977 42901 31980
rect 42935 31977 42947 32011
rect 42889 31971 42947 31977
rect 46934 31968 46940 32020
rect 46992 32008 46998 32020
rect 47029 32011 47087 32017
rect 47029 32008 47041 32011
rect 46992 31980 47041 32008
rect 46992 31968 46998 31980
rect 47029 31977 47041 31980
rect 47075 31977 47087 32011
rect 48682 32008 48688 32020
rect 47029 31971 47087 31977
rect 47688 31980 48688 32008
rect 38565 31943 38623 31949
rect 38565 31909 38577 31943
rect 38611 31940 38623 31943
rect 38838 31940 38844 31952
rect 38611 31912 38844 31940
rect 38611 31909 38623 31912
rect 38565 31903 38623 31909
rect 38838 31900 38844 31912
rect 38896 31900 38902 31952
rect 43070 31940 43076 31952
rect 41984 31912 43076 31940
rect 33778 31872 33784 31884
rect 31036 31844 31156 31872
rect 33060 31844 33784 31872
rect 30469 31807 30527 31813
rect 30469 31773 30481 31807
rect 30515 31773 30527 31807
rect 30469 31767 30527 31773
rect 30653 31807 30711 31813
rect 30653 31773 30665 31807
rect 30699 31804 30711 31807
rect 30699 31776 30972 31804
rect 30699 31773 30711 31776
rect 30653 31767 30711 31773
rect 25308 31739 25366 31745
rect 25308 31705 25320 31739
rect 25354 31736 25366 31739
rect 25498 31736 25504 31748
rect 25354 31708 25504 31736
rect 25354 31705 25366 31708
rect 25308 31699 25366 31705
rect 25498 31696 25504 31708
rect 25556 31696 25562 31748
rect 30944 31668 30972 31776
rect 31036 31736 31064 31844
rect 31113 31807 31171 31813
rect 31113 31773 31125 31807
rect 31159 31804 31171 31807
rect 33060 31804 33088 31844
rect 33778 31832 33784 31844
rect 33836 31872 33842 31884
rect 34698 31872 34704 31884
rect 33836 31844 34704 31872
rect 33836 31832 33842 31844
rect 34698 31832 34704 31844
rect 34756 31832 34762 31884
rect 37182 31872 37188 31884
rect 37143 31844 37188 31872
rect 37182 31832 37188 31844
rect 37240 31832 37246 31884
rect 31159 31776 33088 31804
rect 33137 31807 33195 31813
rect 31159 31773 31171 31776
rect 31113 31767 31171 31773
rect 33137 31773 33149 31807
rect 33183 31773 33195 31807
rect 33137 31767 33195 31773
rect 31358 31739 31416 31745
rect 31358 31736 31370 31739
rect 31036 31708 31370 31736
rect 31358 31705 31370 31708
rect 31404 31705 31416 31739
rect 33152 31736 33180 31767
rect 34514 31764 34520 31816
rect 34572 31804 34578 31816
rect 37458 31813 37464 31816
rect 34957 31807 35015 31813
rect 34957 31804 34969 31807
rect 34572 31776 34969 31804
rect 34572 31764 34578 31776
rect 34957 31773 34969 31776
rect 35003 31773 35015 31807
rect 37452 31804 37464 31813
rect 37419 31776 37464 31804
rect 34957 31767 35015 31773
rect 37452 31767 37464 31776
rect 37458 31764 37464 31767
rect 37516 31764 37522 31816
rect 41984 31813 42012 31912
rect 43070 31900 43076 31912
rect 43128 31900 43134 31952
rect 46750 31900 46756 31952
rect 46808 31940 46814 31952
rect 46808 31912 47532 31940
rect 46808 31900 46814 31912
rect 43533 31875 43591 31881
rect 43533 31872 43545 31875
rect 42168 31844 43545 31872
rect 42168 31813 42196 31844
rect 41969 31807 42027 31813
rect 41969 31773 41981 31807
rect 42015 31773 42027 31807
rect 41969 31767 42027 31773
rect 42153 31807 42211 31813
rect 42153 31773 42165 31807
rect 42199 31773 42211 31807
rect 42153 31767 42211 31773
rect 42242 31764 42248 31816
rect 42300 31804 42306 31816
rect 42812 31813 42840 31844
rect 43533 31841 43545 31844
rect 43579 31841 43591 31875
rect 43533 31835 43591 31841
rect 44361 31875 44419 31881
rect 44361 31841 44373 31875
rect 44407 31872 44419 31875
rect 44407 31844 44588 31872
rect 44407 31841 44419 31844
rect 44361 31835 44419 31841
rect 42797 31807 42855 31813
rect 42300 31776 42345 31804
rect 42300 31764 42306 31776
rect 42797 31773 42809 31807
rect 42843 31773 42855 31807
rect 43438 31804 43444 31816
rect 43399 31776 43444 31804
rect 42797 31767 42855 31773
rect 43438 31764 43444 31776
rect 43496 31764 43502 31816
rect 43622 31804 43628 31816
rect 43583 31776 43628 31804
rect 43622 31764 43628 31776
rect 43680 31764 43686 31816
rect 44266 31804 44272 31816
rect 44227 31776 44272 31804
rect 44266 31764 44272 31776
rect 44324 31764 44330 31816
rect 44450 31804 44456 31816
rect 44411 31776 44456 31804
rect 44450 31764 44456 31776
rect 44508 31764 44514 31816
rect 44560 31804 44588 31844
rect 45186 31832 45192 31884
rect 45244 31872 45250 31884
rect 45281 31875 45339 31881
rect 45281 31872 45293 31875
rect 45244 31844 45293 31872
rect 45244 31832 45250 31844
rect 45281 31841 45293 31844
rect 45327 31841 45339 31875
rect 45281 31835 45339 31841
rect 46658 31832 46664 31884
rect 46716 31872 46722 31884
rect 46716 31844 47440 31872
rect 46716 31832 46722 31844
rect 45002 31804 45008 31816
rect 44560 31776 45008 31804
rect 45002 31764 45008 31776
rect 45060 31804 45066 31816
rect 45465 31807 45523 31813
rect 45465 31804 45477 31807
rect 45060 31776 45477 31804
rect 45060 31764 45066 31776
rect 45465 31773 45477 31776
rect 45511 31773 45523 31807
rect 45465 31767 45523 31773
rect 45649 31807 45707 31813
rect 45649 31773 45661 31807
rect 45695 31804 45707 31807
rect 46750 31804 46756 31816
rect 45695 31776 46756 31804
rect 45695 31773 45707 31776
rect 45649 31767 45707 31773
rect 46750 31764 46756 31776
rect 46808 31764 46814 31816
rect 47412 31813 47440 31844
rect 47504 31813 47532 31912
rect 47213 31807 47271 31813
rect 47213 31773 47225 31807
rect 47259 31804 47271 31807
rect 47397 31807 47455 31813
rect 47259 31776 47348 31804
rect 47259 31773 47271 31776
rect 47213 31767 47271 31773
rect 31358 31699 31416 31705
rect 31726 31708 33180 31736
rect 31726 31668 31754 31708
rect 34698 31696 34704 31748
rect 34756 31736 34762 31748
rect 35802 31736 35808 31748
rect 34756 31708 35808 31736
rect 34756 31696 34762 31708
rect 35802 31696 35808 31708
rect 35860 31696 35866 31748
rect 47320 31736 47348 31776
rect 47397 31773 47409 31807
rect 47443 31773 47455 31807
rect 47397 31767 47455 31773
rect 47489 31807 47547 31813
rect 47489 31773 47501 31807
rect 47535 31773 47547 31807
rect 47688 31804 47716 31980
rect 48682 31968 48688 31980
rect 48740 31968 48746 32020
rect 48866 32008 48872 32020
rect 48827 31980 48872 32008
rect 48866 31968 48872 31980
rect 48924 31968 48930 32020
rect 52273 32011 52331 32017
rect 52273 31977 52285 32011
rect 52319 32008 52331 32011
rect 53098 32008 53104 32020
rect 52319 31980 53104 32008
rect 52319 31977 52331 31980
rect 52273 31971 52331 31977
rect 53098 31968 53104 31980
rect 53156 31968 53162 32020
rect 53558 32008 53564 32020
rect 53519 31980 53564 32008
rect 53558 31968 53564 31980
rect 53616 31968 53622 32020
rect 55398 31968 55404 32020
rect 55456 32008 55462 32020
rect 55456 31980 56180 32008
rect 55456 31968 55462 31980
rect 48133 31943 48191 31949
rect 48133 31909 48145 31943
rect 48179 31940 48191 31943
rect 48314 31940 48320 31952
rect 48179 31912 48320 31940
rect 48179 31909 48191 31912
rect 48133 31903 48191 31909
rect 48314 31900 48320 31912
rect 48372 31940 48378 31952
rect 49418 31940 49424 31952
rect 48372 31912 49424 31940
rect 48372 31900 48378 31912
rect 49418 31900 49424 31912
rect 49476 31900 49482 31952
rect 53193 31943 53251 31949
rect 53193 31909 53205 31943
rect 53239 31940 53251 31943
rect 54754 31940 54760 31952
rect 53239 31912 54760 31940
rect 53239 31909 53251 31912
rect 53193 31903 53251 31909
rect 54754 31900 54760 31912
rect 54812 31900 54818 31952
rect 56042 31900 56048 31952
rect 56100 31900 56106 31952
rect 50617 31875 50675 31881
rect 50617 31841 50629 31875
rect 50663 31872 50675 31875
rect 52733 31875 52791 31881
rect 50663 31844 51074 31872
rect 50663 31841 50675 31844
rect 50617 31835 50675 31841
rect 51046 31816 51074 31844
rect 52733 31841 52745 31875
rect 52779 31872 52791 31875
rect 52822 31872 52828 31884
rect 52779 31844 52828 31872
rect 52779 31841 52791 31844
rect 52733 31835 52791 31841
rect 52822 31832 52828 31844
rect 52880 31832 52886 31884
rect 55677 31875 55735 31881
rect 52932 31844 53696 31872
rect 47946 31804 47952 31816
rect 47489 31767 47547 31773
rect 47596 31776 47716 31804
rect 47907 31776 47952 31804
rect 47596 31736 47624 31776
rect 47946 31764 47952 31776
rect 48004 31764 48010 31816
rect 50890 31804 50896 31816
rect 50851 31776 50896 31804
rect 50890 31764 50896 31776
rect 50948 31764 50954 31816
rect 51046 31776 51080 31816
rect 51074 31764 51080 31776
rect 51132 31764 51138 31816
rect 52457 31807 52515 31813
rect 52457 31773 52469 31807
rect 52503 31804 52515 31807
rect 52546 31804 52552 31816
rect 52503 31776 52552 31804
rect 52503 31773 52515 31776
rect 52457 31767 52515 31773
rect 47320 31708 47624 31736
rect 48777 31739 48835 31745
rect 48777 31705 48789 31739
rect 48823 31736 48835 31739
rect 49970 31736 49976 31748
rect 48823 31708 49976 31736
rect 48823 31705 48835 31708
rect 48777 31699 48835 31705
rect 49970 31696 49976 31708
rect 50028 31696 50034 31748
rect 32490 31668 32496 31680
rect 30944 31640 31754 31668
rect 32451 31640 32496 31668
rect 32490 31628 32496 31640
rect 32548 31628 32554 31680
rect 34974 31628 34980 31680
rect 35032 31668 35038 31680
rect 35710 31668 35716 31680
rect 35032 31640 35716 31668
rect 35032 31628 35038 31640
rect 35710 31628 35716 31640
rect 35768 31628 35774 31680
rect 36081 31671 36139 31677
rect 36081 31637 36093 31671
rect 36127 31668 36139 31671
rect 47118 31668 47124 31680
rect 36127 31640 47124 31668
rect 36127 31637 36139 31640
rect 36081 31631 36139 31637
rect 47118 31628 47124 31640
rect 47176 31628 47182 31680
rect 47302 31628 47308 31680
rect 47360 31668 47366 31680
rect 51350 31668 51356 31680
rect 47360 31640 51356 31668
rect 47360 31628 47366 31640
rect 51350 31628 51356 31640
rect 51408 31668 51414 31680
rect 52472 31668 52500 31767
rect 52546 31764 52552 31776
rect 52604 31764 52610 31816
rect 52638 31764 52644 31816
rect 52696 31804 52702 31816
rect 52932 31804 52960 31844
rect 52696 31776 52960 31804
rect 53377 31807 53435 31813
rect 52696 31764 52702 31776
rect 53377 31773 53389 31807
rect 53423 31804 53435 31807
rect 53466 31804 53472 31816
rect 53423 31776 53472 31804
rect 53423 31773 53435 31776
rect 53377 31767 53435 31773
rect 53466 31764 53472 31776
rect 53524 31764 53530 31816
rect 53668 31813 53696 31844
rect 55677 31841 55689 31875
rect 55723 31872 55735 31875
rect 56060 31872 56088 31900
rect 55723 31844 56088 31872
rect 55723 31841 55735 31844
rect 55677 31835 55735 31841
rect 53653 31807 53711 31813
rect 53653 31773 53665 31807
rect 53699 31804 53711 31807
rect 53742 31804 53748 31816
rect 53699 31776 53748 31804
rect 53699 31773 53711 31776
rect 53653 31767 53711 31773
rect 53742 31764 53748 31776
rect 53800 31764 53806 31816
rect 55858 31804 55864 31816
rect 55819 31776 55864 31804
rect 55858 31764 55864 31776
rect 55916 31764 55922 31816
rect 56045 31807 56103 31813
rect 56045 31773 56057 31807
rect 56091 31804 56103 31807
rect 56152 31804 56180 31980
rect 56091 31776 56180 31804
rect 56091 31773 56103 31776
rect 56045 31767 56103 31773
rect 51408 31640 52500 31668
rect 51408 31628 51414 31640
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 25041 31467 25099 31473
rect 25041 31433 25053 31467
rect 25087 31464 25099 31467
rect 25130 31464 25136 31476
rect 25087 31436 25136 31464
rect 25087 31433 25099 31436
rect 25041 31427 25099 31433
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 28721 31467 28779 31473
rect 28721 31433 28733 31467
rect 28767 31464 28779 31467
rect 28994 31464 29000 31476
rect 28767 31436 29000 31464
rect 28767 31433 28779 31436
rect 28721 31427 28779 31433
rect 28994 31424 29000 31436
rect 29052 31424 29058 31476
rect 30926 31424 30932 31476
rect 30984 31464 30990 31476
rect 32125 31467 32183 31473
rect 32125 31464 32137 31467
rect 30984 31436 32137 31464
rect 30984 31424 30990 31436
rect 32125 31433 32137 31436
rect 32171 31433 32183 31467
rect 35894 31464 35900 31476
rect 32125 31427 32183 31433
rect 35544 31436 35900 31464
rect 26234 31356 26240 31408
rect 26292 31396 26298 31408
rect 28813 31399 28871 31405
rect 28813 31396 28825 31399
rect 26292 31368 28825 31396
rect 26292 31356 26298 31368
rect 28813 31365 28825 31368
rect 28859 31365 28871 31399
rect 31754 31396 31760 31408
rect 28813 31359 28871 31365
rect 30392 31368 31760 31396
rect 25222 31328 25228 31340
rect 25183 31300 25228 31328
rect 25222 31288 25228 31300
rect 25280 31288 25286 31340
rect 27525 31331 27583 31337
rect 27525 31297 27537 31331
rect 27571 31328 27583 31331
rect 27614 31328 27620 31340
rect 27571 31300 27620 31328
rect 27571 31297 27583 31300
rect 27525 31291 27583 31297
rect 27614 31288 27620 31300
rect 27672 31288 27678 31340
rect 27709 31331 27767 31337
rect 27709 31297 27721 31331
rect 27755 31328 27767 31331
rect 28166 31328 28172 31340
rect 27755 31300 28172 31328
rect 27755 31297 27767 31300
rect 27709 31291 27767 31297
rect 28166 31288 28172 31300
rect 28224 31288 28230 31340
rect 30392 31337 30420 31368
rect 31754 31356 31760 31368
rect 31812 31356 31818 31408
rect 31846 31356 31852 31408
rect 31904 31396 31910 31408
rect 32585 31399 32643 31405
rect 32585 31396 32597 31399
rect 31904 31368 32597 31396
rect 31904 31356 31910 31368
rect 32585 31365 32597 31368
rect 32631 31365 32643 31399
rect 32585 31359 32643 31365
rect 30377 31331 30435 31337
rect 30377 31297 30389 31331
rect 30423 31297 30435 31331
rect 30377 31291 30435 31297
rect 31110 31288 31116 31340
rect 31168 31328 31174 31340
rect 31205 31331 31263 31337
rect 31205 31328 31217 31331
rect 31168 31300 31217 31328
rect 31168 31288 31174 31300
rect 31205 31297 31217 31300
rect 31251 31297 31263 31331
rect 31205 31291 31263 31297
rect 31297 31331 31355 31337
rect 31297 31297 31309 31331
rect 31343 31328 31355 31331
rect 32214 31328 32220 31340
rect 31343 31300 32220 31328
rect 31343 31297 31355 31300
rect 31297 31291 31355 31297
rect 32214 31288 32220 31300
rect 32272 31288 32278 31340
rect 32490 31328 32496 31340
rect 32451 31300 32496 31328
rect 32490 31288 32496 31300
rect 32548 31288 32554 31340
rect 34698 31288 34704 31340
rect 34756 31328 34762 31340
rect 34974 31328 34980 31340
rect 34756 31300 34980 31328
rect 34756 31288 34762 31300
rect 34974 31288 34980 31300
rect 35032 31288 35038 31340
rect 35244 31331 35302 31337
rect 35244 31297 35256 31331
rect 35290 31328 35302 31331
rect 35544 31328 35572 31436
rect 35894 31424 35900 31436
rect 35952 31424 35958 31476
rect 39206 31424 39212 31476
rect 39264 31464 39270 31476
rect 39666 31464 39672 31476
rect 39264 31436 39672 31464
rect 39264 31424 39270 31436
rect 39666 31424 39672 31436
rect 39724 31464 39730 31476
rect 39853 31467 39911 31473
rect 39853 31464 39865 31467
rect 39724 31436 39865 31464
rect 39724 31424 39730 31436
rect 39853 31433 39865 31436
rect 39899 31433 39911 31467
rect 39853 31427 39911 31433
rect 40310 31424 40316 31476
rect 40368 31464 40374 31476
rect 40497 31467 40555 31473
rect 40497 31464 40509 31467
rect 40368 31436 40509 31464
rect 40368 31424 40374 31436
rect 40497 31433 40509 31436
rect 40543 31433 40555 31467
rect 40497 31427 40555 31433
rect 43070 31424 43076 31476
rect 43128 31464 43134 31476
rect 43257 31467 43315 31473
rect 43257 31464 43269 31467
rect 43128 31436 43269 31464
rect 43128 31424 43134 31436
rect 43257 31433 43269 31436
rect 43303 31433 43315 31467
rect 43257 31427 43315 31433
rect 43622 31424 43628 31476
rect 43680 31464 43686 31476
rect 45278 31464 45284 31476
rect 43680 31436 45284 31464
rect 43680 31424 43686 31436
rect 37544 31399 37602 31405
rect 37544 31365 37556 31399
rect 37590 31396 37602 31399
rect 37642 31396 37648 31408
rect 37590 31368 37648 31396
rect 37590 31365 37602 31368
rect 37544 31359 37602 31365
rect 37642 31356 37648 31368
rect 37700 31356 37706 31408
rect 41506 31396 41512 31408
rect 39500 31368 41512 31396
rect 35290 31300 35572 31328
rect 35290 31297 35302 31300
rect 35244 31291 35302 31297
rect 35802 31288 35808 31340
rect 35860 31328 35866 31340
rect 37277 31331 37335 31337
rect 37277 31328 37289 31331
rect 35860 31300 37289 31328
rect 35860 31288 35866 31300
rect 37277 31297 37289 31300
rect 37323 31297 37335 31331
rect 37277 31291 37335 31297
rect 38654 31288 38660 31340
rect 38712 31328 38718 31340
rect 39390 31328 39396 31340
rect 38712 31300 39396 31328
rect 38712 31288 38718 31300
rect 39390 31288 39396 31300
rect 39448 31288 39454 31340
rect 39500 31337 39528 31368
rect 41506 31356 41512 31368
rect 41564 31356 41570 31408
rect 39485 31331 39543 31337
rect 39485 31297 39497 31331
rect 39531 31297 39543 31331
rect 39485 31291 39543 31297
rect 39669 31331 39727 31337
rect 39669 31297 39681 31331
rect 39715 31328 39727 31331
rect 40405 31331 40463 31337
rect 40405 31328 40417 31331
rect 39715 31300 40417 31328
rect 39715 31297 39727 31300
rect 39669 31291 39727 31297
rect 40405 31297 40417 31300
rect 40451 31328 40463 31331
rect 40954 31328 40960 31340
rect 40451 31300 40960 31328
rect 40451 31297 40463 31300
rect 40405 31291 40463 31297
rect 28810 31220 28816 31272
rect 28868 31260 28874 31272
rect 28905 31263 28963 31269
rect 28905 31260 28917 31263
rect 28868 31232 28917 31260
rect 28868 31220 28874 31232
rect 28905 31229 28917 31232
rect 28951 31229 28963 31263
rect 28905 31223 28963 31229
rect 30282 31220 30288 31272
rect 30340 31260 30346 31272
rect 31389 31263 31447 31269
rect 31389 31260 31401 31263
rect 30340 31232 31401 31260
rect 30340 31220 30346 31232
rect 31389 31229 31401 31232
rect 31435 31260 31447 31263
rect 32677 31263 32735 31269
rect 31435 31232 32260 31260
rect 31435 31229 31447 31232
rect 31389 31223 31447 31229
rect 32232 31192 32260 31232
rect 32677 31229 32689 31263
rect 32723 31229 32735 31263
rect 32677 31223 32735 31229
rect 32692 31192 32720 31223
rect 32232 31164 32720 31192
rect 38657 31195 38715 31201
rect 38657 31161 38669 31195
rect 38703 31192 38715 31195
rect 39114 31192 39120 31204
rect 38703 31164 39120 31192
rect 38703 31161 38715 31164
rect 38657 31155 38715 31161
rect 39114 31152 39120 31164
rect 39172 31192 39178 31204
rect 39684 31192 39712 31291
rect 40954 31288 40960 31300
rect 41012 31288 41018 31340
rect 43441 31331 43499 31337
rect 43441 31297 43453 31331
rect 43487 31328 43499 31331
rect 43530 31328 43536 31340
rect 43487 31300 43536 31328
rect 43487 31297 43499 31300
rect 43441 31291 43499 31297
rect 43530 31288 43536 31300
rect 43588 31288 43594 31340
rect 43732 31337 43760 31436
rect 45278 31424 45284 31436
rect 45336 31424 45342 31476
rect 46474 31424 46480 31476
rect 46532 31464 46538 31476
rect 46661 31467 46719 31473
rect 46661 31464 46673 31467
rect 46532 31436 46673 31464
rect 46532 31424 46538 31436
rect 46661 31433 46673 31436
rect 46707 31433 46719 31467
rect 48130 31464 48136 31476
rect 48091 31436 48136 31464
rect 46661 31427 46719 31433
rect 48130 31424 48136 31436
rect 48188 31424 48194 31476
rect 49694 31464 49700 31476
rect 49655 31436 49700 31464
rect 49694 31424 49700 31436
rect 49752 31424 49758 31476
rect 50985 31467 51043 31473
rect 50985 31433 50997 31467
rect 51031 31464 51043 31467
rect 51258 31464 51264 31476
rect 51031 31436 51264 31464
rect 51031 31433 51043 31436
rect 50985 31427 51043 31433
rect 51258 31424 51264 31436
rect 51316 31424 51322 31476
rect 51353 31467 51411 31473
rect 51353 31433 51365 31467
rect 51399 31464 51411 31467
rect 53006 31464 53012 31476
rect 51399 31436 53012 31464
rect 51399 31433 51411 31436
rect 51353 31427 51411 31433
rect 49234 31396 49240 31408
rect 44376 31368 49240 31396
rect 44376 31337 44404 31368
rect 49234 31356 49240 31368
rect 49292 31356 49298 31408
rect 50706 31396 50712 31408
rect 50172 31368 50712 31396
rect 43717 31331 43775 31337
rect 43717 31297 43729 31331
rect 43763 31297 43775 31331
rect 43717 31291 43775 31297
rect 44177 31331 44235 31337
rect 44177 31297 44189 31331
rect 44223 31297 44235 31331
rect 44177 31291 44235 31297
rect 44361 31331 44419 31337
rect 44361 31297 44373 31331
rect 44407 31297 44419 31331
rect 44818 31328 44824 31340
rect 44779 31300 44824 31328
rect 44361 31291 44419 31297
rect 44192 31260 44220 31291
rect 44818 31288 44824 31300
rect 44876 31288 44882 31340
rect 46106 31328 46112 31340
rect 46067 31300 46112 31328
rect 46106 31288 46112 31300
rect 46164 31288 46170 31340
rect 47578 31328 47584 31340
rect 47539 31300 47584 31328
rect 47578 31288 47584 31300
rect 47636 31288 47642 31340
rect 47949 31331 48007 31337
rect 47949 31297 47961 31331
rect 47995 31328 48007 31331
rect 48038 31328 48044 31340
rect 47995 31300 48044 31328
rect 47995 31297 48007 31300
rect 47949 31291 48007 31297
rect 44266 31260 44272 31272
rect 44179 31232 44272 31260
rect 44266 31220 44272 31232
rect 44324 31260 44330 31272
rect 44450 31260 44456 31272
rect 44324 31232 44456 31260
rect 44324 31220 44330 31232
rect 44450 31220 44456 31232
rect 44508 31220 44514 31272
rect 45097 31263 45155 31269
rect 45097 31229 45109 31263
rect 45143 31229 45155 31263
rect 45097 31223 45155 31229
rect 39172 31164 39712 31192
rect 39172 31152 39178 31164
rect 43438 31152 43444 31204
rect 43496 31192 43502 31204
rect 43625 31195 43683 31201
rect 43625 31192 43637 31195
rect 43496 31164 43637 31192
rect 43496 31152 43502 31164
rect 43625 31161 43637 31164
rect 43671 31192 43683 31195
rect 45112 31192 45140 31223
rect 45278 31220 45284 31272
rect 45336 31260 45342 31272
rect 46385 31263 46443 31269
rect 46385 31260 46397 31263
rect 45336 31232 46397 31260
rect 45336 31220 45342 31232
rect 46385 31229 46397 31232
rect 46431 31260 46443 31263
rect 47964 31260 47992 31291
rect 48038 31288 48044 31300
rect 48096 31288 48102 31340
rect 49145 31331 49203 31337
rect 49145 31297 49157 31331
rect 49191 31297 49203 31331
rect 49326 31328 49332 31340
rect 49287 31300 49332 31328
rect 49145 31291 49203 31297
rect 46431 31232 47992 31260
rect 49160 31260 49188 31291
rect 49326 31288 49332 31300
rect 49384 31288 49390 31340
rect 49421 31331 49479 31337
rect 49421 31297 49433 31331
rect 49467 31297 49479 31331
rect 49421 31291 49479 31297
rect 49234 31260 49240 31272
rect 49160 31232 49240 31260
rect 46431 31229 46443 31232
rect 46385 31223 46443 31229
rect 49234 31220 49240 31232
rect 49292 31220 49298 31272
rect 49436 31260 49464 31291
rect 49510 31288 49516 31340
rect 49568 31328 49574 31340
rect 50172 31337 50200 31368
rect 50706 31356 50712 31368
rect 50764 31396 50770 31408
rect 51166 31396 51172 31408
rect 50764 31368 51172 31396
rect 50764 31356 50770 31368
rect 51166 31356 51172 31368
rect 51224 31356 51230 31408
rect 51813 31399 51871 31405
rect 51813 31365 51825 31399
rect 51859 31396 51871 31399
rect 51920 31396 51948 31436
rect 53006 31424 53012 31436
rect 53064 31424 53070 31476
rect 53469 31467 53527 31473
rect 53469 31433 53481 31467
rect 53515 31464 53527 31467
rect 54570 31464 54576 31476
rect 53515 31436 54576 31464
rect 53515 31433 53527 31436
rect 53469 31427 53527 31433
rect 54570 31424 54576 31436
rect 54628 31424 54634 31476
rect 55398 31464 55404 31476
rect 54956 31436 55404 31464
rect 51859 31368 51948 31396
rect 51859 31365 51871 31368
rect 51813 31359 51871 31365
rect 52178 31356 52184 31408
rect 52236 31396 52242 31408
rect 52917 31399 52975 31405
rect 52917 31396 52929 31399
rect 52236 31368 52929 31396
rect 52236 31356 52242 31368
rect 52917 31365 52929 31368
rect 52963 31365 52975 31399
rect 53742 31396 53748 31408
rect 53703 31368 53748 31396
rect 52917 31359 52975 31365
rect 53742 31356 53748 31368
rect 53800 31356 53806 31408
rect 50157 31331 50215 31337
rect 49568 31300 49613 31328
rect 49568 31288 49574 31300
rect 50157 31297 50169 31331
rect 50203 31297 50215 31331
rect 50157 31291 50215 31297
rect 50341 31331 50399 31337
rect 50341 31297 50353 31331
rect 50387 31328 50399 31331
rect 50890 31328 50896 31340
rect 50387 31300 50896 31328
rect 50387 31297 50399 31300
rect 50341 31291 50399 31297
rect 50890 31288 50896 31300
rect 50948 31288 50954 31340
rect 51074 31288 51080 31340
rect 51132 31328 51138 31340
rect 51994 31328 52000 31340
rect 51132 31300 51177 31328
rect 51276 31300 51856 31328
rect 51955 31300 52000 31328
rect 51132 31288 51138 31300
rect 49970 31260 49976 31272
rect 49436 31232 49976 31260
rect 49970 31220 49976 31232
rect 50028 31220 50034 31272
rect 50249 31263 50307 31269
rect 50249 31229 50261 31263
rect 50295 31260 50307 31263
rect 51276 31260 51304 31300
rect 50295 31232 51304 31260
rect 51828 31260 51856 31300
rect 51994 31288 52000 31300
rect 52052 31288 52058 31340
rect 52089 31331 52147 31337
rect 52089 31297 52101 31331
rect 52135 31297 52147 31331
rect 52089 31291 52147 31297
rect 52104 31260 52132 31291
rect 52362 31288 52368 31340
rect 52420 31328 52426 31340
rect 52733 31331 52791 31337
rect 52733 31328 52745 31331
rect 52420 31300 52745 31328
rect 52420 31288 52426 31300
rect 52733 31297 52745 31300
rect 52779 31297 52791 31331
rect 52733 31291 52791 31297
rect 53009 31331 53067 31337
rect 53009 31297 53021 31331
rect 53055 31297 53067 31331
rect 53466 31328 53472 31340
rect 53427 31300 53472 31328
rect 53009 31291 53067 31297
rect 51828 31232 52132 31260
rect 50295 31229 50307 31232
rect 50249 31223 50307 31229
rect 49988 31192 50016 31220
rect 50801 31195 50859 31201
rect 50801 31192 50813 31195
rect 43671 31164 46520 31192
rect 49988 31164 50813 31192
rect 43671 31161 43683 31164
rect 43625 31155 43683 31161
rect 27706 31084 27712 31136
rect 27764 31124 27770 31136
rect 27893 31127 27951 31133
rect 27893 31124 27905 31127
rect 27764 31096 27905 31124
rect 27764 31084 27770 31096
rect 27893 31093 27905 31096
rect 27939 31093 27951 31127
rect 27893 31087 27951 31093
rect 28353 31127 28411 31133
rect 28353 31093 28365 31127
rect 28399 31124 28411 31127
rect 28994 31124 29000 31136
rect 28399 31096 29000 31124
rect 28399 31093 28411 31096
rect 28353 31087 28411 31093
rect 28994 31084 29000 31096
rect 29052 31084 29058 31136
rect 30190 31124 30196 31136
rect 30151 31096 30196 31124
rect 30190 31084 30196 31096
rect 30248 31084 30254 31136
rect 30837 31127 30895 31133
rect 30837 31093 30849 31127
rect 30883 31124 30895 31127
rect 32306 31124 32312 31136
rect 30883 31096 32312 31124
rect 30883 31093 30895 31096
rect 30837 31087 30895 31093
rect 32306 31084 32312 31096
rect 32364 31084 32370 31136
rect 36357 31127 36415 31133
rect 36357 31093 36369 31127
rect 36403 31124 36415 31127
rect 36630 31124 36636 31136
rect 36403 31096 36636 31124
rect 36403 31093 36415 31096
rect 36357 31087 36415 31093
rect 36630 31084 36636 31096
rect 36688 31084 36694 31136
rect 38838 31084 38844 31136
rect 38896 31124 38902 31136
rect 39022 31124 39028 31136
rect 38896 31096 39028 31124
rect 38896 31084 38902 31096
rect 39022 31084 39028 31096
rect 39080 31124 39086 31136
rect 39482 31124 39488 31136
rect 39080 31096 39488 31124
rect 39080 31084 39086 31096
rect 39482 31084 39488 31096
rect 39540 31084 39546 31136
rect 44174 31124 44180 31136
rect 44135 31096 44180 31124
rect 44174 31084 44180 31096
rect 44232 31084 44238 31136
rect 44358 31084 44364 31136
rect 44416 31124 44422 31136
rect 44726 31124 44732 31136
rect 44416 31096 44732 31124
rect 44416 31084 44422 31096
rect 44726 31084 44732 31096
rect 44784 31084 44790 31136
rect 46492 31133 46520 31164
rect 50801 31161 50813 31164
rect 50847 31161 50859 31195
rect 50801 31155 50859 31161
rect 51813 31195 51871 31201
rect 51813 31161 51825 31195
rect 51859 31192 51871 31195
rect 51902 31192 51908 31204
rect 51859 31164 51908 31192
rect 51859 31161 51871 31164
rect 51813 31155 51871 31161
rect 51902 31152 51908 31164
rect 51960 31152 51966 31204
rect 52733 31195 52791 31201
rect 52733 31161 52745 31195
rect 52779 31192 52791 31195
rect 52822 31192 52828 31204
rect 52779 31164 52828 31192
rect 52779 31161 52791 31164
rect 52733 31155 52791 31161
rect 52822 31152 52828 31164
rect 52880 31152 52886 31204
rect 46477 31127 46535 31133
rect 46477 31093 46489 31127
rect 46523 31124 46535 31127
rect 47949 31127 48007 31133
rect 47949 31124 47961 31127
rect 46523 31096 47961 31124
rect 46523 31093 46535 31096
rect 46477 31087 46535 31093
rect 47949 31093 47961 31096
rect 47995 31124 48007 31127
rect 48222 31124 48228 31136
rect 47995 31096 48228 31124
rect 47995 31093 48007 31096
rect 47949 31087 48007 31093
rect 48222 31084 48228 31096
rect 48280 31084 48286 31136
rect 51166 31084 51172 31136
rect 51224 31124 51230 31136
rect 53024 31124 53052 31291
rect 53466 31288 53472 31300
rect 53524 31288 53530 31340
rect 53558 31288 53564 31340
rect 53616 31328 53622 31340
rect 54956 31337 54984 31436
rect 55398 31424 55404 31436
rect 55456 31424 55462 31476
rect 55582 31464 55588 31476
rect 55543 31436 55588 31464
rect 55582 31424 55588 31436
rect 55640 31424 55646 31476
rect 55953 31467 56011 31473
rect 55953 31433 55965 31467
rect 55999 31464 56011 31467
rect 56134 31464 56140 31476
rect 55999 31436 56140 31464
rect 55999 31433 56011 31436
rect 55953 31427 56011 31433
rect 56134 31424 56140 31436
rect 56192 31424 56198 31476
rect 56594 31464 56600 31476
rect 56555 31436 56600 31464
rect 56594 31424 56600 31436
rect 56652 31424 56658 31476
rect 55033 31399 55091 31405
rect 55033 31365 55045 31399
rect 55079 31396 55091 31399
rect 55858 31396 55864 31408
rect 55079 31368 55864 31396
rect 55079 31365 55091 31368
rect 55033 31359 55091 31365
rect 55858 31356 55864 31368
rect 55916 31356 55922 31408
rect 56689 31399 56747 31405
rect 56689 31396 56701 31399
rect 56060 31368 56701 31396
rect 56060 31340 56088 31368
rect 56689 31365 56701 31368
rect 56735 31365 56747 31399
rect 56689 31359 56747 31365
rect 54941 31331 54999 31337
rect 53616 31300 53661 31328
rect 53616 31288 53622 31300
rect 54941 31297 54953 31331
rect 54987 31297 54999 31331
rect 54941 31291 54999 31297
rect 55125 31331 55183 31337
rect 55125 31297 55137 31331
rect 55171 31297 55183 31331
rect 55766 31328 55772 31340
rect 55727 31300 55772 31328
rect 55125 31291 55183 31297
rect 53650 31152 53656 31204
rect 53708 31192 53714 31204
rect 55140 31192 55168 31291
rect 55766 31288 55772 31300
rect 55824 31288 55830 31340
rect 56042 31288 56048 31340
rect 56100 31328 56106 31340
rect 56505 31331 56563 31337
rect 56100 31300 56145 31328
rect 56100 31288 56106 31300
rect 56505 31297 56517 31331
rect 56551 31297 56563 31331
rect 56505 31291 56563 31297
rect 56781 31331 56839 31337
rect 56781 31297 56793 31331
rect 56827 31297 56839 31331
rect 56781 31291 56839 31297
rect 55784 31260 55812 31288
rect 56520 31260 56548 31291
rect 55784 31232 56548 31260
rect 55582 31192 55588 31204
rect 53708 31164 55588 31192
rect 53708 31152 53714 31164
rect 55582 31152 55588 31164
rect 55640 31152 55646 31204
rect 56134 31152 56140 31204
rect 56192 31192 56198 31204
rect 56796 31192 56824 31291
rect 56192 31164 56824 31192
rect 56192 31152 56198 31164
rect 51224 31096 53052 31124
rect 51224 31084 51230 31096
rect 56318 31084 56324 31136
rect 56376 31124 56382 31136
rect 58069 31127 58127 31133
rect 58069 31124 58081 31127
rect 56376 31096 58081 31124
rect 56376 31084 56382 31096
rect 58069 31093 58081 31096
rect 58115 31093 58127 31127
rect 58069 31087 58127 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 28166 30880 28172 30932
rect 28224 30920 28230 30932
rect 28261 30923 28319 30929
rect 28261 30920 28273 30923
rect 28224 30892 28273 30920
rect 28224 30880 28230 30892
rect 28261 30889 28273 30892
rect 28307 30889 28319 30923
rect 28261 30883 28319 30889
rect 31202 30880 31208 30932
rect 31260 30920 31266 30932
rect 32401 30923 32459 30929
rect 32401 30920 32413 30923
rect 31260 30892 32413 30920
rect 31260 30880 31266 30892
rect 32401 30889 32413 30892
rect 32447 30889 32459 30923
rect 36722 30920 36728 30932
rect 36683 30892 36728 30920
rect 32401 30883 32459 30889
rect 36722 30880 36728 30892
rect 36780 30880 36786 30932
rect 39022 30920 39028 30932
rect 38983 30892 39028 30920
rect 39022 30880 39028 30892
rect 39080 30880 39086 30932
rect 44269 30923 44327 30929
rect 44269 30889 44281 30923
rect 44315 30920 44327 30923
rect 44818 30920 44824 30932
rect 44315 30892 44824 30920
rect 44315 30889 44327 30892
rect 44269 30883 44327 30889
rect 44818 30880 44824 30892
rect 44876 30880 44882 30932
rect 46290 30920 46296 30932
rect 46251 30892 46296 30920
rect 46290 30880 46296 30892
rect 46348 30880 46354 30932
rect 47946 30880 47952 30932
rect 48004 30920 48010 30932
rect 48225 30923 48283 30929
rect 48225 30920 48237 30923
rect 48004 30892 48237 30920
rect 48004 30880 48010 30892
rect 48225 30889 48237 30892
rect 48271 30889 48283 30923
rect 49142 30920 49148 30932
rect 49103 30892 49148 30920
rect 48225 30883 48283 30889
rect 49142 30880 49148 30892
rect 49200 30880 49206 30932
rect 50706 30920 50712 30932
rect 50667 30892 50712 30920
rect 50706 30880 50712 30892
rect 50764 30880 50770 30932
rect 51350 30920 51356 30932
rect 51311 30892 51356 30920
rect 51350 30880 51356 30892
rect 51408 30880 51414 30932
rect 52273 30923 52331 30929
rect 52273 30889 52285 30923
rect 52319 30889 52331 30923
rect 52273 30883 52331 30889
rect 52457 30923 52515 30929
rect 52457 30889 52469 30923
rect 52503 30920 52515 30923
rect 52638 30920 52644 30932
rect 52503 30892 52644 30920
rect 52503 30889 52515 30892
rect 52457 30883 52515 30889
rect 39390 30852 39396 30864
rect 38948 30824 39396 30852
rect 38948 30796 38976 30824
rect 39390 30812 39396 30824
rect 39448 30812 39454 30864
rect 41322 30812 41328 30864
rect 41380 30852 41386 30864
rect 48774 30852 48780 30864
rect 41380 30824 48780 30852
rect 41380 30812 41386 30824
rect 48774 30812 48780 30824
rect 48832 30852 48838 30864
rect 49007 30855 49065 30861
rect 49007 30852 49019 30855
rect 48832 30824 49019 30852
rect 48832 30812 48838 30824
rect 49007 30821 49019 30824
rect 49053 30821 49065 30855
rect 49007 30815 49065 30821
rect 28905 30787 28963 30793
rect 28905 30753 28917 30787
rect 28951 30784 28963 30787
rect 30282 30784 30288 30796
rect 28951 30756 30288 30784
rect 28951 30753 28963 30756
rect 28905 30747 28963 30753
rect 30282 30744 30288 30756
rect 30340 30744 30346 30796
rect 38930 30784 38936 30796
rect 38891 30756 38936 30784
rect 38930 30744 38936 30756
rect 38988 30744 38994 30796
rect 40221 30787 40279 30793
rect 40221 30784 40233 30787
rect 39040 30756 40233 30784
rect 27706 30716 27712 30728
rect 27667 30688 27712 30716
rect 27706 30676 27712 30688
rect 27764 30676 27770 30728
rect 28721 30719 28779 30725
rect 28721 30685 28733 30719
rect 28767 30716 28779 30719
rect 29270 30716 29276 30728
rect 28767 30688 29276 30716
rect 28767 30685 28779 30688
rect 28721 30679 28779 30685
rect 29270 30676 29276 30688
rect 29328 30676 29334 30728
rect 31021 30719 31079 30725
rect 31021 30685 31033 30719
rect 31067 30716 31079 30719
rect 34698 30716 34704 30728
rect 31067 30688 34704 30716
rect 31067 30685 31079 30688
rect 31021 30679 31079 30685
rect 34698 30676 34704 30688
rect 34756 30676 34762 30728
rect 35526 30676 35532 30728
rect 35584 30716 35590 30728
rect 35713 30719 35771 30725
rect 35713 30716 35725 30719
rect 35584 30688 35725 30716
rect 35584 30676 35590 30688
rect 35713 30685 35725 30688
rect 35759 30685 35771 30719
rect 36630 30716 36636 30728
rect 36591 30688 36636 30716
rect 35713 30679 35771 30685
rect 36630 30676 36636 30688
rect 36688 30676 36694 30728
rect 36722 30676 36728 30728
rect 36780 30716 36786 30728
rect 37553 30719 37611 30725
rect 37553 30716 37565 30719
rect 36780 30688 37565 30716
rect 36780 30676 36786 30688
rect 37553 30685 37565 30688
rect 37599 30685 37611 30719
rect 37553 30679 37611 30685
rect 38841 30719 38899 30725
rect 38841 30685 38853 30719
rect 38887 30716 38899 30719
rect 39040 30716 39068 30756
rect 40221 30753 40233 30756
rect 40267 30784 40279 30787
rect 41506 30784 41512 30796
rect 40267 30756 41512 30784
rect 40267 30753 40279 30756
rect 40221 30747 40279 30753
rect 41506 30744 41512 30756
rect 41564 30744 41570 30796
rect 44542 30784 44548 30796
rect 43640 30756 44548 30784
rect 38887 30688 39068 30716
rect 38887 30685 38899 30688
rect 38841 30679 38899 30685
rect 39114 30676 39120 30728
rect 39172 30716 39178 30728
rect 39172 30688 39217 30716
rect 39172 30676 39178 30688
rect 39298 30676 39304 30728
rect 39356 30716 39362 30728
rect 39942 30716 39948 30728
rect 39356 30688 39948 30716
rect 39356 30676 39362 30688
rect 39942 30676 39948 30688
rect 40000 30676 40006 30728
rect 41233 30719 41291 30725
rect 41233 30685 41245 30719
rect 41279 30685 41291 30719
rect 43438 30716 43444 30728
rect 43399 30688 43444 30716
rect 41233 30679 41291 30685
rect 30190 30608 30196 30660
rect 30248 30648 30254 30660
rect 31266 30651 31324 30657
rect 31266 30648 31278 30651
rect 30248 30620 31278 30648
rect 30248 30608 30254 30620
rect 31266 30617 31278 30620
rect 31312 30617 31324 30651
rect 31266 30611 31324 30617
rect 35989 30651 36047 30657
rect 35989 30617 36001 30651
rect 36035 30648 36047 30651
rect 37182 30648 37188 30660
rect 36035 30620 37188 30648
rect 36035 30617 36047 30620
rect 35989 30611 36047 30617
rect 37182 30608 37188 30620
rect 37240 30608 37246 30660
rect 40402 30648 40408 30660
rect 37752 30620 40408 30648
rect 27522 30580 27528 30592
rect 27483 30552 27528 30580
rect 27522 30540 27528 30552
rect 27580 30540 27586 30592
rect 28350 30540 28356 30592
rect 28408 30580 28414 30592
rect 28629 30583 28687 30589
rect 28629 30580 28641 30583
rect 28408 30552 28641 30580
rect 28408 30540 28414 30552
rect 28629 30549 28641 30552
rect 28675 30549 28687 30583
rect 37090 30580 37096 30592
rect 37051 30552 37096 30580
rect 28629 30543 28687 30549
rect 37090 30540 37096 30552
rect 37148 30540 37154 30592
rect 37752 30589 37780 30620
rect 40402 30608 40408 30620
rect 40460 30648 40466 30660
rect 41248 30648 41276 30679
rect 43438 30676 43444 30688
rect 43496 30676 43502 30728
rect 43640 30725 43668 30756
rect 44542 30744 44548 30756
rect 44600 30744 44606 30796
rect 45278 30784 45284 30796
rect 45239 30756 45284 30784
rect 45278 30744 45284 30756
rect 45336 30744 45342 30796
rect 51074 30784 51080 30796
rect 48148 30756 51080 30784
rect 43625 30719 43683 30725
rect 43625 30685 43637 30719
rect 43671 30685 43683 30719
rect 43625 30679 43683 30685
rect 44085 30719 44143 30725
rect 44085 30685 44097 30719
rect 44131 30685 44143 30719
rect 44266 30716 44272 30728
rect 44227 30688 44272 30716
rect 44085 30679 44143 30685
rect 40460 30620 41276 30648
rect 44100 30648 44128 30679
rect 44266 30676 44272 30688
rect 44324 30716 44330 30728
rect 45005 30719 45063 30725
rect 45005 30716 45017 30719
rect 44324 30688 45017 30716
rect 44324 30676 44330 30688
rect 45005 30685 45017 30688
rect 45051 30685 45063 30719
rect 46474 30716 46480 30728
rect 46435 30688 46480 30716
rect 45005 30679 45063 30685
rect 46474 30676 46480 30688
rect 46532 30676 46538 30728
rect 46750 30716 46756 30728
rect 46711 30688 46756 30716
rect 46750 30676 46756 30688
rect 46808 30676 46814 30728
rect 47118 30676 47124 30728
rect 47176 30716 47182 30728
rect 48148 30725 48176 30756
rect 51074 30744 51080 30756
rect 51132 30784 51138 30796
rect 51132 30756 51488 30784
rect 51132 30744 51138 30756
rect 48133 30719 48191 30725
rect 48133 30716 48145 30719
rect 47176 30688 48145 30716
rect 47176 30676 47182 30688
rect 48133 30685 48145 30688
rect 48179 30685 48191 30719
rect 48866 30716 48872 30728
rect 48827 30688 48872 30716
rect 48133 30679 48191 30685
rect 48866 30676 48872 30688
rect 48924 30676 48930 30728
rect 49329 30719 49387 30725
rect 49329 30685 49341 30719
rect 49375 30716 49387 30719
rect 49694 30716 49700 30728
rect 49375 30688 49700 30716
rect 49375 30685 49387 30688
rect 49329 30679 49387 30685
rect 49694 30676 49700 30688
rect 49752 30676 49758 30728
rect 51166 30676 51172 30728
rect 51224 30716 51230 30728
rect 51460 30725 51488 30756
rect 51261 30719 51319 30725
rect 51261 30716 51273 30719
rect 51224 30688 51273 30716
rect 51224 30676 51230 30688
rect 51261 30685 51273 30688
rect 51307 30685 51319 30719
rect 51261 30679 51319 30685
rect 51445 30719 51503 30725
rect 51445 30685 51457 30719
rect 51491 30685 51503 30719
rect 52288 30716 52316 30883
rect 52638 30880 52644 30892
rect 52696 30880 52702 30932
rect 55769 30923 55827 30929
rect 55769 30889 55781 30923
rect 55815 30920 55827 30923
rect 56042 30920 56048 30932
rect 55815 30892 56048 30920
rect 55815 30889 55827 30892
rect 55769 30883 55827 30889
rect 56042 30880 56048 30892
rect 56100 30880 56106 30932
rect 56318 30784 56324 30796
rect 56279 30756 56324 30784
rect 56318 30744 56324 30756
rect 56376 30744 56382 30796
rect 51445 30679 51503 30685
rect 51552 30688 52316 30716
rect 54481 30719 54539 30725
rect 44358 30648 44364 30660
rect 44100 30620 44364 30648
rect 40460 30608 40466 30620
rect 44358 30608 44364 30620
rect 44416 30608 44422 30660
rect 44726 30648 44732 30660
rect 44468 30620 44732 30648
rect 37737 30583 37795 30589
rect 37737 30549 37749 30583
rect 37783 30549 37795 30583
rect 37737 30543 37795 30549
rect 39301 30583 39359 30589
rect 39301 30549 39313 30583
rect 39347 30580 39359 30583
rect 40218 30580 40224 30592
rect 39347 30552 40224 30580
rect 39347 30549 39359 30552
rect 39301 30543 39359 30549
rect 40218 30540 40224 30552
rect 40276 30540 40282 30592
rect 40586 30540 40592 30592
rect 40644 30580 40650 30592
rect 41322 30580 41328 30592
rect 40644 30552 41328 30580
rect 40644 30540 40650 30552
rect 41322 30540 41328 30552
rect 41380 30540 41386 30592
rect 43530 30580 43536 30592
rect 43491 30552 43536 30580
rect 43530 30540 43536 30552
rect 43588 30540 43594 30592
rect 44468 30589 44496 30620
rect 44726 30608 44732 30620
rect 44784 30608 44790 30660
rect 47762 30608 47768 30660
rect 47820 30648 47826 30660
rect 48884 30648 48912 30676
rect 47820 30620 48912 30648
rect 50617 30651 50675 30657
rect 47820 30608 47826 30620
rect 50617 30617 50629 30651
rect 50663 30648 50675 30651
rect 50982 30648 50988 30660
rect 50663 30620 50988 30648
rect 50663 30617 50675 30620
rect 50617 30611 50675 30617
rect 50982 30608 50988 30620
rect 51040 30648 51046 30660
rect 51552 30648 51580 30688
rect 54481 30685 54493 30719
rect 54527 30685 54539 30719
rect 54662 30716 54668 30728
rect 54623 30688 54668 30716
rect 54481 30679 54539 30685
rect 52086 30648 52092 30660
rect 51040 30620 51580 30648
rect 52047 30620 52092 30648
rect 51040 30608 51046 30620
rect 52086 30608 52092 30620
rect 52144 30608 52150 30660
rect 52362 30657 52368 30660
rect 52305 30651 52368 30657
rect 52305 30617 52317 30651
rect 52351 30617 52368 30651
rect 52305 30611 52368 30617
rect 52362 30608 52368 30611
rect 52420 30608 52426 30660
rect 54496 30648 54524 30679
rect 54662 30676 54668 30688
rect 54720 30676 54726 30728
rect 55582 30716 55588 30728
rect 55543 30688 55588 30716
rect 55582 30676 55588 30688
rect 55640 30676 55646 30728
rect 54754 30648 54760 30660
rect 54496 30620 54760 30648
rect 54754 30608 54760 30620
rect 54812 30608 54818 30660
rect 55398 30648 55404 30660
rect 55359 30620 55404 30648
rect 55398 30608 55404 30620
rect 55456 30608 55462 30660
rect 56505 30651 56563 30657
rect 56505 30617 56517 30651
rect 56551 30648 56563 30651
rect 57974 30648 57980 30660
rect 56551 30620 57980 30648
rect 56551 30617 56563 30620
rect 56505 30611 56563 30617
rect 57974 30608 57980 30620
rect 58032 30608 58038 30660
rect 58158 30648 58164 30660
rect 58119 30620 58164 30648
rect 58158 30608 58164 30620
rect 58216 30608 58222 30660
rect 44453 30583 44511 30589
rect 44453 30549 44465 30583
rect 44499 30549 44511 30583
rect 44453 30543 44511 30549
rect 46566 30540 46572 30592
rect 46624 30580 46630 30592
rect 46661 30583 46719 30589
rect 46661 30580 46673 30583
rect 46624 30552 46673 30580
rect 46624 30540 46630 30552
rect 46661 30549 46673 30552
rect 46707 30549 46719 30583
rect 46661 30543 46719 30549
rect 49329 30583 49387 30589
rect 49329 30549 49341 30583
rect 49375 30580 49387 30583
rect 50154 30580 50160 30592
rect 49375 30552 50160 30580
rect 49375 30549 49387 30552
rect 49329 30543 49387 30549
rect 50154 30540 50160 30552
rect 50212 30540 50218 30592
rect 54202 30540 54208 30592
rect 54260 30580 54266 30592
rect 54573 30583 54631 30589
rect 54573 30580 54585 30583
rect 54260 30552 54585 30580
rect 54260 30540 54266 30552
rect 54573 30549 54585 30552
rect 54619 30549 54631 30583
rect 54573 30543 54631 30549
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 28350 30376 28356 30388
rect 28311 30348 28356 30376
rect 28350 30336 28356 30348
rect 28408 30336 28414 30388
rect 35526 30336 35532 30388
rect 35584 30376 35590 30388
rect 38654 30376 38660 30388
rect 35584 30348 36676 30376
rect 38615 30348 38660 30376
rect 35584 30336 35590 30348
rect 27240 30311 27298 30317
rect 27240 30277 27252 30311
rect 27286 30308 27298 30311
rect 27522 30308 27528 30320
rect 27286 30280 27528 30308
rect 27286 30277 27298 30280
rect 27240 30271 27298 30277
rect 27522 30268 27528 30280
rect 27580 30268 27586 30320
rect 34146 30317 34152 30320
rect 34140 30271 34152 30317
rect 34204 30308 34210 30320
rect 36648 30317 36676 30348
rect 38654 30336 38660 30348
rect 38712 30376 38718 30388
rect 38838 30376 38844 30388
rect 38712 30348 38844 30376
rect 38712 30336 38718 30348
rect 38838 30336 38844 30348
rect 38896 30376 38902 30388
rect 40310 30376 40316 30388
rect 38896 30348 38976 30376
rect 40271 30348 40316 30376
rect 38896 30336 38902 30348
rect 36633 30311 36691 30317
rect 34204 30280 34240 30308
rect 34146 30268 34152 30271
rect 34204 30268 34210 30280
rect 36633 30277 36645 30311
rect 36679 30277 36691 30311
rect 37090 30308 37096 30320
rect 36633 30271 36691 30277
rect 36740 30280 37096 30308
rect 2406 30240 2412 30252
rect 2367 30212 2412 30240
rect 2406 30200 2412 30212
rect 2464 30200 2470 30252
rect 24578 30200 24584 30252
rect 24636 30240 24642 30252
rect 25961 30243 26019 30249
rect 25961 30240 25973 30243
rect 24636 30212 25973 30240
rect 24636 30200 24642 30212
rect 25961 30209 25973 30212
rect 26007 30209 26019 30243
rect 26970 30240 26976 30252
rect 26931 30212 26976 30240
rect 25961 30203 26019 30209
rect 26970 30200 26976 30212
rect 27028 30200 27034 30252
rect 28074 30200 28080 30252
rect 28132 30240 28138 30252
rect 28810 30240 28816 30252
rect 28132 30212 28816 30240
rect 28132 30200 28138 30212
rect 28810 30200 28816 30212
rect 28868 30240 28874 30252
rect 28997 30243 29055 30249
rect 28997 30240 29009 30243
rect 28868 30212 29009 30240
rect 28868 30200 28874 30212
rect 28997 30209 29009 30212
rect 29043 30209 29055 30243
rect 28997 30203 29055 30209
rect 30837 30243 30895 30249
rect 30837 30209 30849 30243
rect 30883 30240 30895 30243
rect 30883 30212 31754 30240
rect 30883 30209 30895 30212
rect 30837 30203 30895 30209
rect 30852 30172 30880 30203
rect 31110 30172 31116 30184
rect 28920 30144 30880 30172
rect 31071 30144 31116 30172
rect 1946 30036 1952 30048
rect 1907 30008 1952 30036
rect 1946 29996 1952 30008
rect 2004 29996 2010 30048
rect 2130 29996 2136 30048
rect 2188 30036 2194 30048
rect 2501 30039 2559 30045
rect 2501 30036 2513 30039
rect 2188 30008 2513 30036
rect 2188 29996 2194 30008
rect 2501 30005 2513 30008
rect 2547 30005 2559 30039
rect 26050 30036 26056 30048
rect 26011 30008 26056 30036
rect 2501 29999 2559 30005
rect 26050 29996 26056 30008
rect 26108 29996 26114 30048
rect 26421 30039 26479 30045
rect 26421 30005 26433 30039
rect 26467 30036 26479 30039
rect 28920 30036 28948 30144
rect 31110 30132 31116 30144
rect 31168 30132 31174 30184
rect 31726 30172 31754 30212
rect 33778 30200 33784 30252
rect 33836 30240 33842 30252
rect 36740 30249 36768 30280
rect 37090 30268 37096 30280
rect 37148 30308 37154 30320
rect 37148 30280 38884 30308
rect 37148 30268 37154 30280
rect 33873 30243 33931 30249
rect 33873 30240 33885 30243
rect 33836 30212 33885 30240
rect 33836 30200 33842 30212
rect 33873 30209 33885 30212
rect 33919 30209 33931 30243
rect 33873 30203 33931 30209
rect 36449 30243 36507 30249
rect 36449 30209 36461 30243
rect 36495 30209 36507 30243
rect 36449 30203 36507 30209
rect 36725 30243 36783 30249
rect 36725 30209 36737 30243
rect 36771 30209 36783 30243
rect 36725 30203 36783 30209
rect 37553 30243 37611 30249
rect 37553 30209 37565 30243
rect 37599 30209 37611 30243
rect 37553 30203 37611 30209
rect 38381 30243 38439 30249
rect 38381 30209 38393 30243
rect 38427 30240 38439 30243
rect 38654 30240 38660 30252
rect 38427 30212 38660 30240
rect 38427 30209 38439 30212
rect 38381 30203 38439 30209
rect 31938 30172 31944 30184
rect 31726 30144 31944 30172
rect 31938 30132 31944 30144
rect 31996 30132 32002 30184
rect 36464 30172 36492 30203
rect 37568 30172 37596 30203
rect 38654 30200 38660 30212
rect 38712 30200 38718 30252
rect 38856 30249 38884 30280
rect 38841 30243 38899 30249
rect 38841 30209 38853 30243
rect 38887 30209 38899 30243
rect 38948 30240 38976 30348
rect 40310 30336 40316 30348
rect 40368 30336 40374 30388
rect 43438 30336 43444 30388
rect 43496 30376 43502 30388
rect 44542 30376 44548 30388
rect 43496 30348 44312 30376
rect 43496 30336 43502 30348
rect 41874 30308 41880 30320
rect 41835 30280 41880 30308
rect 41874 30268 41880 30280
rect 41932 30268 41938 30320
rect 43257 30311 43315 30317
rect 43257 30277 43269 30311
rect 43303 30308 43315 30311
rect 43530 30308 43536 30320
rect 43303 30280 43536 30308
rect 43303 30277 43315 30280
rect 43257 30271 43315 30277
rect 43530 30268 43536 30280
rect 43588 30268 43594 30320
rect 39301 30243 39359 30249
rect 39301 30240 39313 30243
rect 38948 30212 39313 30240
rect 38841 30203 38899 30209
rect 39301 30209 39313 30212
rect 39347 30209 39359 30243
rect 39942 30240 39948 30252
rect 39903 30212 39948 30240
rect 39301 30203 39359 30209
rect 39942 30200 39948 30212
rect 40000 30200 40006 30252
rect 41509 30243 41567 30249
rect 41509 30209 41521 30243
rect 41555 30209 41567 30243
rect 41509 30203 41567 30209
rect 36464 30144 37596 30172
rect 30653 30107 30711 30113
rect 30653 30073 30665 30107
rect 30699 30104 30711 30107
rect 31662 30104 31668 30116
rect 30699 30076 31668 30104
rect 30699 30073 30711 30076
rect 30653 30067 30711 30073
rect 31662 30064 31668 30076
rect 31720 30064 31726 30116
rect 37568 30104 37596 30144
rect 38473 30175 38531 30181
rect 38473 30141 38485 30175
rect 38519 30172 38531 30175
rect 38562 30172 38568 30184
rect 38519 30144 38568 30172
rect 38519 30141 38531 30144
rect 38473 30135 38531 30141
rect 38562 30132 38568 30144
rect 38620 30132 38626 30184
rect 38749 30175 38807 30181
rect 38749 30141 38761 30175
rect 38795 30172 38807 30175
rect 38795 30144 39528 30172
rect 38795 30141 38807 30144
rect 38749 30135 38807 30141
rect 39393 30107 39451 30113
rect 39393 30104 39405 30107
rect 37568 30076 39405 30104
rect 39393 30073 39405 30076
rect 39439 30073 39451 30107
rect 39500 30104 39528 30144
rect 40494 30132 40500 30184
rect 40552 30172 40558 30184
rect 40552 30144 41414 30172
rect 40552 30132 40558 30144
rect 39500 30076 40540 30104
rect 39393 30067 39451 30073
rect 40512 30048 40540 30076
rect 29086 30036 29092 30048
rect 26467 30008 28948 30036
rect 29047 30008 29092 30036
rect 26467 30005 26479 30008
rect 26421 29999 26479 30005
rect 29086 29996 29092 30008
rect 29144 29996 29150 30048
rect 29457 30039 29515 30045
rect 29457 30005 29469 30039
rect 29503 30036 29515 30039
rect 30466 30036 30472 30048
rect 29503 30008 30472 30036
rect 29503 30005 29515 30008
rect 29457 29999 29515 30005
rect 30466 29996 30472 30008
rect 30524 29996 30530 30048
rect 30834 29996 30840 30048
rect 30892 30036 30898 30048
rect 31021 30039 31079 30045
rect 31021 30036 31033 30039
rect 30892 30008 31033 30036
rect 30892 29996 30898 30008
rect 31021 30005 31033 30008
rect 31067 30005 31079 30039
rect 31021 29999 31079 30005
rect 35253 30039 35311 30045
rect 35253 30005 35265 30039
rect 35299 30036 35311 30039
rect 35802 30036 35808 30048
rect 35299 30008 35808 30036
rect 35299 30005 35311 30008
rect 35253 29999 35311 30005
rect 35802 29996 35808 30008
rect 35860 29996 35866 30048
rect 36446 30036 36452 30048
rect 36407 30008 36452 30036
rect 36446 29996 36452 30008
rect 36504 29996 36510 30048
rect 37642 30036 37648 30048
rect 37603 30008 37648 30036
rect 37642 29996 37648 30008
rect 37700 29996 37706 30048
rect 37734 29996 37740 30048
rect 37792 30036 37798 30048
rect 38197 30039 38255 30045
rect 38197 30036 38209 30039
rect 37792 30008 38209 30036
rect 37792 29996 37798 30008
rect 38197 30005 38209 30008
rect 38243 30005 38255 30039
rect 40310 30036 40316 30048
rect 40271 30008 40316 30036
rect 38197 29999 38255 30005
rect 40310 29996 40316 30008
rect 40368 29996 40374 30048
rect 40494 30036 40500 30048
rect 40455 30008 40500 30036
rect 40494 29996 40500 30008
rect 40552 29996 40558 30048
rect 41386 30036 41414 30144
rect 41524 30104 41552 30203
rect 41598 30200 41604 30252
rect 41656 30240 41662 30252
rect 41693 30243 41751 30249
rect 41693 30240 41705 30243
rect 41656 30212 41705 30240
rect 41656 30200 41662 30212
rect 41693 30209 41705 30212
rect 41739 30209 41751 30243
rect 42426 30240 42432 30252
rect 42387 30212 42432 30240
rect 41693 30203 41751 30209
rect 42426 30200 42432 30212
rect 42484 30200 42490 30252
rect 42521 30243 42579 30249
rect 42521 30209 42533 30243
rect 42567 30240 42579 30243
rect 42702 30240 42708 30252
rect 42567 30212 42708 30240
rect 42567 30209 42579 30212
rect 42521 30203 42579 30209
rect 42702 30200 42708 30212
rect 42760 30200 42766 30252
rect 42797 30243 42855 30249
rect 42797 30209 42809 30243
rect 42843 30240 42855 30243
rect 43441 30243 43499 30249
rect 43441 30240 43453 30243
rect 42843 30212 43453 30240
rect 42843 30209 42855 30212
rect 42797 30203 42855 30209
rect 43441 30209 43453 30212
rect 43487 30240 43499 30243
rect 43990 30240 43996 30252
rect 43487 30212 43996 30240
rect 43487 30209 43499 30212
rect 43441 30203 43499 30209
rect 43990 30200 43996 30212
rect 44048 30200 44054 30252
rect 44177 30243 44235 30249
rect 44177 30209 44189 30243
rect 44223 30209 44235 30243
rect 44284 30240 44312 30348
rect 44376 30348 44548 30376
rect 44376 30317 44404 30348
rect 44542 30336 44548 30348
rect 44600 30376 44606 30388
rect 45462 30376 45468 30388
rect 44600 30348 45468 30376
rect 44600 30336 44606 30348
rect 45462 30336 45468 30348
rect 45520 30336 45526 30388
rect 49142 30336 49148 30388
rect 49200 30376 49206 30388
rect 49513 30379 49571 30385
rect 49513 30376 49525 30379
rect 49200 30348 49525 30376
rect 49200 30336 49206 30348
rect 49513 30345 49525 30348
rect 49559 30345 49571 30379
rect 55766 30376 55772 30388
rect 55727 30348 55772 30376
rect 49513 30339 49571 30345
rect 55766 30336 55772 30348
rect 55824 30336 55830 30388
rect 44361 30311 44419 30317
rect 44361 30277 44373 30311
rect 44407 30277 44419 30311
rect 44361 30271 44419 30277
rect 44821 30311 44879 30317
rect 44821 30277 44833 30311
rect 44867 30308 44879 30311
rect 44910 30308 44916 30320
rect 44867 30280 44916 30308
rect 44867 30277 44879 30280
rect 44821 30271 44879 30277
rect 44910 30268 44916 30280
rect 44968 30268 44974 30320
rect 48961 30311 49019 30317
rect 48961 30277 48973 30311
rect 49007 30308 49019 30311
rect 49326 30308 49332 30320
rect 49007 30280 49332 30308
rect 49007 30277 49019 30280
rect 48961 30271 49019 30277
rect 49326 30268 49332 30280
rect 49384 30268 49390 30320
rect 50982 30308 50988 30320
rect 49436 30280 50988 30308
rect 45005 30243 45063 30249
rect 44284 30212 44956 30240
rect 44177 30203 44235 30209
rect 42058 30132 42064 30184
rect 42116 30172 42122 30184
rect 42613 30175 42671 30181
rect 42613 30172 42625 30175
rect 42116 30144 42625 30172
rect 42116 30132 42122 30144
rect 42613 30141 42625 30144
rect 42659 30172 42671 30175
rect 43346 30172 43352 30184
rect 42659 30144 43352 30172
rect 42659 30141 42671 30144
rect 42613 30135 42671 30141
rect 43346 30132 43352 30144
rect 43404 30172 43410 30184
rect 43625 30175 43683 30181
rect 43625 30172 43637 30175
rect 43404 30144 43637 30172
rect 43404 30132 43410 30144
rect 43625 30141 43637 30144
rect 43671 30172 43683 30175
rect 43806 30172 43812 30184
rect 43671 30144 43812 30172
rect 43671 30141 43683 30144
rect 43625 30135 43683 30141
rect 43806 30132 43812 30144
rect 43864 30132 43870 30184
rect 42797 30107 42855 30113
rect 42797 30104 42809 30107
rect 41524 30076 42809 30104
rect 42797 30073 42809 30076
rect 42843 30073 42855 30107
rect 42797 30067 42855 30073
rect 43530 30064 43536 30116
rect 43588 30104 43594 30116
rect 44192 30104 44220 30203
rect 44928 30184 44956 30212
rect 45005 30209 45017 30243
rect 45051 30209 45063 30243
rect 45186 30240 45192 30252
rect 45147 30212 45192 30240
rect 45005 30203 45063 30209
rect 44910 30132 44916 30184
rect 44968 30132 44974 30184
rect 45020 30172 45048 30203
rect 45186 30200 45192 30212
rect 45244 30200 45250 30252
rect 45281 30243 45339 30249
rect 45281 30209 45293 30243
rect 45327 30240 45339 30243
rect 46750 30240 46756 30252
rect 45327 30212 46756 30240
rect 45327 30209 45339 30212
rect 45281 30203 45339 30209
rect 46750 30200 46756 30212
rect 46808 30200 46814 30252
rect 47946 30200 47952 30252
rect 48004 30240 48010 30252
rect 48041 30243 48099 30249
rect 48041 30240 48053 30243
rect 48004 30212 48053 30240
rect 48004 30200 48010 30212
rect 48041 30209 48053 30212
rect 48087 30209 48099 30243
rect 48041 30203 48099 30209
rect 48225 30243 48283 30249
rect 48225 30209 48237 30243
rect 48271 30209 48283 30243
rect 48225 30203 48283 30209
rect 45094 30172 45100 30184
rect 45020 30144 45100 30172
rect 45094 30132 45100 30144
rect 45152 30132 45158 30184
rect 48240 30172 48268 30203
rect 48682 30200 48688 30252
rect 48740 30240 48746 30252
rect 48777 30243 48835 30249
rect 48777 30240 48789 30243
rect 48740 30212 48789 30240
rect 48740 30200 48746 30212
rect 48777 30209 48789 30212
rect 48823 30209 48835 30243
rect 48777 30203 48835 30209
rect 49234 30200 49240 30252
rect 49292 30240 49298 30252
rect 49436 30249 49464 30280
rect 50982 30268 50988 30280
rect 51040 30268 51046 30320
rect 54202 30268 54208 30320
rect 54260 30308 54266 30320
rect 55585 30311 55643 30317
rect 55585 30308 55597 30311
rect 54260 30280 55597 30308
rect 54260 30268 54266 30280
rect 55585 30277 55597 30280
rect 55631 30277 55643 30311
rect 57974 30308 57980 30320
rect 57935 30280 57980 30308
rect 55585 30271 55643 30277
rect 57974 30268 57980 30280
rect 58032 30268 58038 30320
rect 49421 30243 49479 30249
rect 49421 30240 49433 30243
rect 49292 30212 49433 30240
rect 49292 30200 49298 30212
rect 49421 30209 49433 30212
rect 49467 30209 49479 30243
rect 49421 30203 49479 30209
rect 49510 30200 49516 30252
rect 49568 30240 49574 30252
rect 49605 30243 49663 30249
rect 49605 30240 49617 30243
rect 49568 30212 49617 30240
rect 49568 30200 49574 30212
rect 49605 30209 49617 30212
rect 49651 30209 49663 30243
rect 49605 30203 49663 30209
rect 51077 30243 51135 30249
rect 51077 30209 51089 30243
rect 51123 30240 51135 30243
rect 51258 30240 51264 30252
rect 51123 30212 51264 30240
rect 51123 30209 51135 30212
rect 51077 30203 51135 30209
rect 51258 30200 51264 30212
rect 51316 30240 51322 30252
rect 52086 30240 52092 30252
rect 51316 30212 52092 30240
rect 51316 30200 51322 30212
rect 52086 30200 52092 30212
rect 52144 30200 52150 30252
rect 54662 30240 54668 30252
rect 54623 30212 54668 30240
rect 54662 30200 54668 30212
rect 54720 30200 54726 30252
rect 54754 30200 54760 30252
rect 54812 30240 54818 30252
rect 54941 30243 54999 30249
rect 54812 30212 54857 30240
rect 54812 30200 54818 30212
rect 54941 30209 54953 30243
rect 54987 30240 54999 30243
rect 55401 30243 55459 30249
rect 55401 30240 55413 30243
rect 54987 30212 55413 30240
rect 54987 30209 54999 30212
rect 54941 30203 54999 30209
rect 55401 30209 55413 30212
rect 55447 30209 55459 30243
rect 55401 30203 55459 30209
rect 56686 30200 56692 30252
rect 56744 30240 56750 30252
rect 57149 30243 57207 30249
rect 57149 30240 57161 30243
rect 56744 30212 57161 30240
rect 56744 30200 56750 30212
rect 57149 30209 57161 30212
rect 57195 30240 57207 30243
rect 57330 30240 57336 30252
rect 57195 30212 57336 30240
rect 57195 30209 57207 30212
rect 57149 30203 57207 30209
rect 57330 30200 57336 30212
rect 57388 30200 57394 30252
rect 57606 30200 57612 30252
rect 57664 30240 57670 30252
rect 57885 30243 57943 30249
rect 57885 30240 57897 30243
rect 57664 30212 57897 30240
rect 57664 30200 57670 30212
rect 57885 30209 57897 30212
rect 57931 30209 57943 30243
rect 57885 30203 57943 30209
rect 49970 30172 49976 30184
rect 48240 30144 49976 30172
rect 49970 30132 49976 30144
rect 50028 30132 50034 30184
rect 50798 30172 50804 30184
rect 50759 30144 50804 30172
rect 50798 30132 50804 30144
rect 50856 30132 50862 30184
rect 49510 30104 49516 30116
rect 43588 30076 44220 30104
rect 47964 30076 49516 30104
rect 43588 30064 43594 30076
rect 47964 30036 47992 30076
rect 49510 30064 49516 30076
rect 49568 30064 49574 30116
rect 49602 30064 49608 30116
rect 49660 30104 49666 30116
rect 51994 30104 52000 30116
rect 49660 30076 52000 30104
rect 49660 30064 49666 30076
rect 51994 30064 52000 30076
rect 52052 30064 52058 30116
rect 48130 30036 48136 30048
rect 41386 30008 47992 30036
rect 48091 30008 48136 30036
rect 48130 29996 48136 30008
rect 48188 29996 48194 30048
rect 56502 29996 56508 30048
rect 56560 30036 56566 30048
rect 57241 30039 57299 30045
rect 57241 30036 57253 30039
rect 56560 30008 57253 30036
rect 56560 29996 56566 30008
rect 57241 30005 57253 30008
rect 57287 30005 57299 30039
rect 57241 29999 57299 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 31113 29835 31171 29841
rect 31113 29801 31125 29835
rect 31159 29832 31171 29835
rect 31846 29832 31852 29844
rect 31159 29804 31852 29832
rect 31159 29801 31171 29804
rect 31113 29795 31171 29801
rect 31846 29792 31852 29804
rect 31904 29792 31910 29844
rect 38565 29835 38623 29841
rect 38565 29801 38577 29835
rect 38611 29832 38623 29835
rect 38654 29832 38660 29844
rect 38611 29804 38660 29832
rect 38611 29801 38623 29804
rect 38565 29795 38623 29801
rect 38654 29792 38660 29804
rect 38712 29792 38718 29844
rect 38746 29792 38752 29844
rect 38804 29832 38810 29844
rect 39758 29832 39764 29844
rect 38804 29804 39764 29832
rect 38804 29792 38810 29804
rect 39758 29792 39764 29804
rect 39816 29792 39822 29844
rect 42242 29792 42248 29844
rect 42300 29832 42306 29844
rect 42429 29835 42487 29841
rect 42429 29832 42441 29835
rect 42300 29804 42441 29832
rect 42300 29792 42306 29804
rect 42429 29801 42441 29804
rect 42475 29801 42487 29835
rect 42429 29795 42487 29801
rect 43441 29835 43499 29841
rect 43441 29801 43453 29835
rect 43487 29832 43499 29835
rect 45186 29832 45192 29844
rect 43487 29804 45192 29832
rect 43487 29801 43499 29804
rect 43441 29795 43499 29801
rect 45186 29792 45192 29804
rect 45244 29832 45250 29844
rect 45244 29804 46336 29832
rect 45244 29792 45250 29804
rect 26896 29736 28120 29764
rect 24578 29588 24584 29640
rect 24636 29628 24642 29640
rect 26896 29637 26924 29736
rect 28092 29708 28120 29736
rect 30834 29724 30840 29776
rect 30892 29764 30898 29776
rect 31757 29767 31815 29773
rect 31757 29764 31769 29767
rect 30892 29736 31769 29764
rect 30892 29724 30898 29736
rect 31757 29733 31769 29736
rect 31803 29733 31815 29767
rect 31757 29727 31815 29733
rect 36446 29724 36452 29776
rect 36504 29764 36510 29776
rect 40034 29764 40040 29776
rect 36504 29736 40040 29764
rect 36504 29724 36510 29736
rect 40034 29724 40040 29736
rect 40092 29724 40098 29776
rect 40218 29764 40224 29776
rect 40179 29736 40224 29764
rect 40218 29724 40224 29736
rect 40276 29724 40282 29776
rect 40402 29724 40408 29776
rect 40460 29764 40466 29776
rect 40460 29736 43484 29764
rect 40460 29724 40466 29736
rect 43456 29708 43484 29736
rect 43530 29724 43536 29776
rect 43588 29764 43594 29776
rect 43588 29736 45232 29764
rect 43588 29724 43594 29736
rect 27982 29696 27988 29708
rect 27943 29668 27988 29696
rect 27982 29656 27988 29668
rect 28040 29656 28046 29708
rect 28074 29656 28080 29708
rect 28132 29696 28138 29708
rect 28132 29668 28225 29696
rect 28132 29656 28138 29668
rect 31110 29656 31116 29708
rect 31168 29696 31174 29708
rect 31938 29696 31944 29708
rect 31168 29668 31708 29696
rect 31899 29668 31944 29696
rect 31168 29656 31174 29668
rect 26881 29631 26939 29637
rect 26881 29628 26893 29631
rect 24636 29600 26893 29628
rect 24636 29588 24642 29600
rect 26881 29597 26893 29600
rect 26927 29597 26939 29631
rect 26881 29591 26939 29597
rect 27893 29631 27951 29637
rect 27893 29597 27905 29631
rect 27939 29628 27951 29631
rect 28350 29628 28356 29640
rect 27939 29600 28356 29628
rect 27939 29597 27951 29600
rect 27893 29591 27951 29597
rect 28350 29588 28356 29600
rect 28408 29588 28414 29640
rect 30834 29628 30840 29640
rect 29840 29600 30840 29628
rect 27065 29563 27123 29569
rect 27065 29529 27077 29563
rect 27111 29560 27123 29563
rect 27338 29560 27344 29572
rect 27111 29532 27344 29560
rect 27111 29529 27123 29532
rect 27065 29523 27123 29529
rect 27338 29520 27344 29532
rect 27396 29560 27402 29572
rect 29840 29560 29868 29600
rect 30834 29588 30840 29600
rect 30892 29588 30898 29640
rect 31680 29637 31708 29668
rect 31938 29656 31944 29668
rect 31996 29656 32002 29708
rect 36630 29696 36636 29708
rect 36096 29668 36636 29696
rect 31021 29631 31079 29637
rect 31021 29597 31033 29631
rect 31067 29628 31079 29631
rect 31665 29631 31723 29637
rect 31067 29600 31340 29628
rect 31067 29597 31079 29600
rect 31021 29591 31079 29597
rect 27396 29532 29868 29560
rect 27396 29520 27402 29532
rect 30466 29520 30472 29572
rect 30524 29560 30530 29572
rect 31205 29563 31263 29569
rect 31205 29560 31217 29563
rect 30524 29532 31217 29560
rect 30524 29520 30530 29532
rect 31205 29529 31217 29532
rect 31251 29529 31263 29563
rect 31312 29560 31340 29600
rect 31665 29597 31677 29631
rect 31711 29597 31723 29631
rect 31665 29591 31723 29597
rect 33134 29588 33140 29640
rect 33192 29628 33198 29640
rect 36096 29637 36124 29668
rect 36630 29656 36636 29668
rect 36688 29696 36694 29708
rect 36725 29699 36783 29705
rect 36725 29696 36737 29699
rect 36688 29668 36737 29696
rect 36688 29656 36694 29668
rect 36725 29665 36737 29668
rect 36771 29665 36783 29699
rect 36725 29659 36783 29665
rect 38470 29656 38476 29708
rect 38528 29696 38534 29708
rect 39209 29699 39267 29705
rect 39209 29696 39221 29699
rect 38528 29668 39221 29696
rect 38528 29656 38534 29668
rect 39209 29665 39221 29668
rect 39255 29696 39267 29699
rect 40494 29696 40500 29708
rect 39255 29668 40500 29696
rect 39255 29665 39267 29668
rect 39209 29659 39267 29665
rect 40494 29656 40500 29668
rect 40552 29656 40558 29708
rect 42153 29699 42211 29705
rect 42153 29665 42165 29699
rect 42199 29696 42211 29699
rect 42610 29696 42616 29708
rect 42199 29668 42616 29696
rect 42199 29665 42211 29668
rect 42153 29659 42211 29665
rect 42610 29656 42616 29668
rect 42668 29656 42674 29708
rect 43438 29656 43444 29708
rect 43496 29656 43502 29708
rect 45097 29699 45155 29705
rect 45097 29696 45109 29699
rect 44008 29668 45109 29696
rect 44008 29640 44036 29668
rect 45097 29665 45109 29668
rect 45143 29665 45155 29699
rect 45097 29659 45155 29665
rect 33597 29631 33655 29637
rect 33597 29628 33609 29631
rect 33192 29600 33609 29628
rect 33192 29588 33198 29600
rect 33597 29597 33609 29600
rect 33643 29597 33655 29631
rect 33597 29591 33655 29597
rect 36081 29631 36139 29637
rect 36081 29597 36093 29631
rect 36127 29597 36139 29631
rect 36998 29628 37004 29640
rect 36959 29600 37004 29628
rect 36081 29591 36139 29597
rect 36998 29588 37004 29600
rect 37056 29588 37062 29640
rect 37182 29588 37188 29640
rect 37240 29628 37246 29640
rect 38746 29628 38752 29640
rect 37240 29600 38752 29628
rect 37240 29588 37246 29600
rect 38746 29588 38752 29600
rect 38804 29588 38810 29640
rect 38841 29631 38899 29637
rect 38841 29597 38853 29631
rect 38887 29597 38899 29631
rect 40037 29631 40095 29637
rect 40037 29628 40049 29631
rect 38841 29591 38899 29597
rect 38948 29600 40049 29628
rect 31754 29560 31760 29572
rect 31312 29532 31760 29560
rect 31205 29523 31263 29529
rect 31754 29520 31760 29532
rect 31812 29560 31818 29572
rect 32490 29560 32496 29572
rect 31812 29532 32496 29560
rect 31812 29520 31818 29532
rect 32490 29520 32496 29532
rect 32548 29520 32554 29572
rect 33686 29560 33692 29572
rect 33647 29532 33692 29560
rect 33686 29520 33692 29532
rect 33744 29520 33750 29572
rect 37016 29560 37044 29588
rect 38856 29560 38884 29591
rect 37016 29532 38884 29560
rect 27525 29495 27583 29501
rect 27525 29461 27537 29495
rect 27571 29492 27583 29495
rect 28534 29492 28540 29504
rect 27571 29464 28540 29492
rect 27571 29461 27583 29464
rect 27525 29455 27583 29461
rect 28534 29452 28540 29464
rect 28592 29452 28598 29504
rect 31938 29492 31944 29504
rect 31899 29464 31944 29492
rect 31938 29452 31944 29464
rect 31996 29452 32002 29504
rect 36173 29495 36231 29501
rect 36173 29461 36185 29495
rect 36219 29492 36231 29495
rect 36262 29492 36268 29504
rect 36219 29464 36268 29492
rect 36219 29461 36231 29464
rect 36173 29455 36231 29461
rect 36262 29452 36268 29464
rect 36320 29492 36326 29504
rect 38948 29492 38976 29600
rect 40037 29597 40049 29600
rect 40083 29597 40095 29631
rect 40037 29591 40095 29597
rect 39574 29560 39580 29572
rect 39040 29532 39580 29560
rect 39040 29501 39068 29532
rect 39574 29520 39580 29532
rect 39632 29520 39638 29572
rect 40052 29560 40080 29591
rect 40126 29588 40132 29640
rect 40184 29628 40190 29640
rect 40313 29631 40371 29637
rect 40184 29600 40229 29628
rect 40184 29588 40190 29600
rect 40313 29597 40325 29631
rect 40359 29628 40371 29631
rect 40402 29628 40408 29640
rect 40359 29600 40408 29628
rect 40359 29597 40371 29600
rect 40313 29591 40371 29597
rect 40402 29588 40408 29600
rect 40460 29588 40466 29640
rect 40954 29628 40960 29640
rect 40915 29600 40960 29628
rect 40954 29588 40960 29600
rect 41012 29588 41018 29640
rect 42058 29628 42064 29640
rect 42019 29600 42064 29628
rect 42058 29588 42064 29600
rect 42116 29588 42122 29640
rect 43626 29628 43684 29631
rect 43806 29628 43812 29640
rect 43569 29625 43684 29628
rect 43569 29600 43638 29625
rect 40218 29560 40224 29572
rect 40052 29532 40224 29560
rect 40218 29520 40224 29532
rect 40276 29520 40282 29572
rect 43162 29520 43168 29572
rect 43220 29560 43226 29572
rect 43569 29560 43597 29600
rect 43626 29591 43638 29600
rect 43672 29591 43684 29625
rect 43767 29600 43812 29628
rect 43626 29585 43684 29591
rect 43806 29588 43812 29600
rect 43864 29588 43870 29640
rect 43990 29628 43996 29640
rect 43951 29600 43996 29628
rect 43990 29588 43996 29600
rect 44048 29588 44054 29640
rect 44085 29631 44143 29637
rect 44085 29597 44097 29631
rect 44131 29628 44143 29631
rect 44174 29628 44180 29640
rect 44131 29600 44180 29628
rect 44131 29597 44143 29600
rect 44085 29591 44143 29597
rect 44174 29588 44180 29600
rect 44232 29588 44238 29640
rect 44910 29588 44916 29640
rect 44968 29628 44974 29640
rect 45204 29637 45232 29736
rect 45005 29631 45063 29637
rect 45005 29628 45017 29631
rect 44968 29600 45017 29628
rect 44968 29588 44974 29600
rect 45005 29597 45017 29600
rect 45051 29597 45063 29631
rect 45005 29591 45063 29597
rect 45189 29631 45247 29637
rect 45189 29597 45201 29631
rect 45235 29597 45247 29631
rect 45189 29591 45247 29597
rect 43220 29532 43597 29560
rect 43220 29520 43226 29532
rect 43714 29520 43720 29572
rect 43772 29560 43778 29572
rect 46308 29560 46336 29804
rect 46382 29792 46388 29844
rect 46440 29832 46446 29844
rect 46937 29835 46995 29841
rect 46937 29832 46949 29835
rect 46440 29804 46949 29832
rect 46440 29792 46446 29804
rect 46937 29801 46949 29804
rect 46983 29801 46995 29835
rect 46937 29795 46995 29801
rect 47578 29792 47584 29844
rect 47636 29832 47642 29844
rect 47949 29835 48007 29841
rect 47949 29832 47961 29835
rect 47636 29804 47961 29832
rect 47636 29792 47642 29804
rect 47949 29801 47961 29804
rect 47995 29801 48007 29835
rect 47949 29795 48007 29801
rect 52089 29835 52147 29841
rect 52089 29801 52101 29835
rect 52135 29832 52147 29835
rect 52730 29832 52736 29844
rect 52135 29804 52736 29832
rect 52135 29801 52147 29804
rect 52089 29795 52147 29801
rect 52730 29792 52736 29804
rect 52788 29792 52794 29844
rect 54018 29832 54024 29844
rect 53979 29804 54024 29832
rect 54018 29792 54024 29804
rect 54076 29792 54082 29844
rect 55398 29832 55404 29844
rect 55359 29804 55404 29832
rect 55398 29792 55404 29804
rect 55456 29792 55462 29844
rect 46750 29764 46756 29776
rect 46400 29736 46756 29764
rect 46400 29637 46428 29736
rect 46750 29724 46756 29736
rect 46808 29724 46814 29776
rect 47854 29764 47860 29776
rect 47596 29736 47860 29764
rect 47596 29696 47624 29736
rect 47854 29724 47860 29736
rect 47912 29724 47918 29776
rect 50154 29724 50160 29776
rect 50212 29764 50218 29776
rect 50212 29736 52776 29764
rect 50212 29724 50218 29736
rect 46768 29668 47624 29696
rect 47673 29699 47731 29705
rect 46768 29637 46796 29668
rect 47673 29665 47685 29699
rect 47719 29696 47731 29699
rect 48774 29696 48780 29708
rect 47719 29668 48780 29696
rect 47719 29665 47731 29668
rect 47673 29659 47731 29665
rect 48774 29656 48780 29668
rect 48832 29656 48838 29708
rect 52748 29705 52776 29736
rect 51353 29699 51411 29705
rect 51353 29665 51365 29699
rect 51399 29696 51411 29699
rect 52733 29699 52791 29705
rect 51399 29668 52132 29696
rect 51399 29665 51411 29668
rect 51353 29659 51411 29665
rect 46385 29631 46443 29637
rect 46385 29597 46397 29631
rect 46431 29597 46443 29631
rect 46385 29591 46443 29597
rect 46753 29631 46811 29637
rect 46753 29597 46765 29631
rect 46799 29597 46811 29631
rect 47578 29628 47584 29640
rect 47491 29600 47584 29628
rect 46753 29591 46811 29597
rect 47578 29588 47584 29600
rect 47636 29628 47642 29640
rect 48130 29628 48136 29640
rect 47636 29600 48136 29628
rect 47636 29588 47642 29600
rect 48130 29588 48136 29600
rect 48188 29588 48194 29640
rect 51166 29588 51172 29640
rect 51224 29628 51230 29640
rect 51261 29631 51319 29637
rect 51261 29628 51273 29631
rect 51224 29600 51273 29628
rect 51224 29588 51230 29600
rect 51261 29597 51273 29600
rect 51307 29597 51319 29631
rect 51442 29628 51448 29640
rect 51403 29600 51448 29628
rect 51261 29591 51319 29597
rect 51442 29588 51448 29600
rect 51500 29588 51506 29640
rect 51905 29631 51963 29637
rect 51905 29597 51917 29631
rect 51951 29597 51963 29631
rect 52104 29628 52132 29668
rect 52733 29665 52745 29699
rect 52779 29665 52791 29699
rect 52733 29659 52791 29665
rect 53193 29699 53251 29705
rect 53193 29665 53205 29699
rect 53239 29696 53251 29699
rect 54018 29696 54024 29708
rect 53239 29668 54024 29696
rect 53239 29665 53251 29668
rect 53193 29659 53251 29665
rect 54018 29656 54024 29668
rect 54076 29696 54082 29708
rect 56502 29696 56508 29708
rect 54076 29668 54524 29696
rect 56463 29668 56508 29696
rect 54076 29656 54082 29668
rect 52825 29631 52883 29637
rect 52825 29628 52837 29631
rect 52104 29600 52837 29628
rect 51905 29591 51963 29597
rect 52825 29597 52837 29600
rect 52871 29597 52883 29631
rect 54202 29628 54208 29640
rect 54163 29600 54208 29628
rect 52825 29591 52883 29597
rect 46566 29560 46572 29572
rect 43772 29532 43817 29560
rect 46308 29532 46572 29560
rect 43772 29520 43778 29532
rect 46566 29520 46572 29532
rect 46624 29520 46630 29572
rect 46661 29563 46719 29569
rect 46661 29529 46673 29563
rect 46707 29560 46719 29563
rect 47762 29560 47768 29572
rect 46707 29532 47768 29560
rect 46707 29529 46719 29532
rect 46661 29523 46719 29529
rect 47762 29520 47768 29532
rect 47820 29520 47826 29572
rect 51920 29560 51948 29591
rect 54202 29588 54208 29600
rect 54260 29588 54266 29640
rect 54496 29637 54524 29668
rect 56502 29656 56508 29668
rect 56560 29656 56566 29708
rect 57882 29696 57888 29708
rect 57843 29668 57888 29696
rect 57882 29656 57888 29668
rect 57940 29656 57946 29708
rect 54481 29631 54539 29637
rect 54481 29597 54493 29631
rect 54527 29597 54539 29631
rect 55306 29628 55312 29640
rect 55267 29600 55312 29628
rect 54481 29591 54539 29597
rect 55306 29588 55312 29600
rect 55364 29588 55370 29640
rect 55490 29628 55496 29640
rect 55451 29600 55496 29628
rect 55490 29588 55496 29600
rect 55548 29628 55554 29640
rect 56134 29628 56140 29640
rect 55548 29600 56140 29628
rect 55548 29588 55554 29600
rect 56134 29588 56140 29600
rect 56192 29588 56198 29640
rect 56318 29628 56324 29640
rect 56279 29600 56324 29628
rect 56318 29588 56324 29600
rect 56376 29588 56382 29640
rect 52454 29560 52460 29572
rect 51920 29532 52460 29560
rect 52454 29520 52460 29532
rect 52512 29520 52518 29572
rect 36320 29464 38976 29492
rect 39025 29495 39083 29501
rect 36320 29452 36326 29464
rect 39025 29461 39037 29495
rect 39071 29461 39083 29495
rect 39025 29455 39083 29461
rect 39117 29495 39175 29501
rect 39117 29461 39129 29495
rect 39163 29492 39175 29495
rect 39206 29492 39212 29504
rect 39163 29464 39212 29492
rect 39163 29461 39175 29464
rect 39117 29455 39175 29461
rect 39206 29452 39212 29464
rect 39264 29452 39270 29504
rect 39298 29452 39304 29504
rect 39356 29492 39362 29504
rect 39853 29495 39911 29501
rect 39853 29492 39865 29495
rect 39356 29464 39865 29492
rect 39356 29452 39362 29464
rect 39853 29461 39865 29464
rect 39899 29461 39911 29495
rect 41046 29492 41052 29504
rect 41007 29464 41052 29492
rect 39853 29455 39911 29461
rect 41046 29452 41052 29464
rect 41104 29492 41110 29504
rect 43530 29492 43536 29504
rect 41104 29464 43536 29492
rect 41104 29452 41110 29464
rect 43530 29452 43536 29464
rect 43588 29452 43594 29504
rect 49878 29452 49884 29504
rect 49936 29492 49942 29504
rect 53006 29492 53012 29504
rect 49936 29464 53012 29492
rect 49936 29452 49942 29464
rect 53006 29452 53012 29464
rect 53064 29452 53070 29504
rect 54386 29492 54392 29504
rect 54347 29464 54392 29492
rect 54386 29452 54392 29464
rect 54444 29452 54450 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 28074 29248 28080 29300
rect 28132 29288 28138 29300
rect 28353 29291 28411 29297
rect 28353 29288 28365 29291
rect 28132 29260 28365 29288
rect 28132 29248 28138 29260
rect 28353 29257 28365 29260
rect 28399 29257 28411 29291
rect 28353 29251 28411 29257
rect 32493 29291 32551 29297
rect 32493 29257 32505 29291
rect 32539 29288 32551 29291
rect 42610 29288 42616 29300
rect 32539 29260 33364 29288
rect 32539 29257 32551 29260
rect 32493 29251 32551 29257
rect 2130 29220 2136 29232
rect 2091 29192 2136 29220
rect 2130 29180 2136 29192
rect 2188 29180 2194 29232
rect 33336 29229 33364 29260
rect 38672 29260 39620 29288
rect 42571 29260 42616 29288
rect 33321 29223 33379 29229
rect 33321 29189 33333 29223
rect 33367 29189 33379 29223
rect 33321 29183 33379 29189
rect 38565 29223 38623 29229
rect 38565 29189 38577 29223
rect 38611 29220 38623 29223
rect 38672 29220 38700 29260
rect 38611 29192 38700 29220
rect 38611 29189 38623 29192
rect 38565 29183 38623 29189
rect 1946 29152 1952 29164
rect 1907 29124 1952 29152
rect 1946 29112 1952 29124
rect 2004 29112 2010 29164
rect 24578 29152 24584 29164
rect 24539 29124 24584 29152
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 26970 29152 26976 29164
rect 26931 29124 26976 29152
rect 26970 29112 26976 29124
rect 27028 29112 27034 29164
rect 27246 29161 27252 29164
rect 27240 29115 27252 29161
rect 27304 29152 27310 29164
rect 27304 29124 27340 29152
rect 27246 29112 27252 29115
rect 27304 29112 27310 29124
rect 30466 29112 30472 29164
rect 30524 29152 30530 29164
rect 30837 29155 30895 29161
rect 30837 29152 30849 29155
rect 30524 29124 30849 29152
rect 30524 29112 30530 29124
rect 30837 29121 30849 29124
rect 30883 29121 30895 29155
rect 30837 29115 30895 29121
rect 31018 29112 31024 29164
rect 31076 29152 31082 29164
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31076 29124 32137 29152
rect 31076 29112 31082 29124
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 37277 29155 37335 29161
rect 37277 29121 37289 29155
rect 37323 29152 37335 29155
rect 37918 29152 37924 29164
rect 37323 29124 37924 29152
rect 37323 29121 37335 29124
rect 37277 29115 37335 29121
rect 37918 29112 37924 29124
rect 37976 29112 37982 29164
rect 38470 29152 38476 29164
rect 38431 29124 38476 29152
rect 38470 29112 38476 29124
rect 38528 29112 38534 29164
rect 38657 29155 38715 29161
rect 38657 29152 38669 29155
rect 38580 29124 38669 29152
rect 2774 29084 2780 29096
rect 2735 29056 2780 29084
rect 2774 29044 2780 29056
rect 2832 29044 2838 29096
rect 24765 29087 24823 29093
rect 24765 29053 24777 29087
rect 24811 29084 24823 29087
rect 25222 29084 25228 29096
rect 24811 29056 25228 29084
rect 24811 29053 24823 29056
rect 24765 29047 24823 29053
rect 25222 29044 25228 29056
rect 25280 29044 25286 29096
rect 25317 29087 25375 29093
rect 25317 29053 25329 29087
rect 25363 29053 25375 29087
rect 25317 29047 25375 29053
rect 31113 29087 31171 29093
rect 31113 29053 31125 29087
rect 31159 29084 31171 29087
rect 31754 29084 31760 29096
rect 31159 29056 31760 29084
rect 31159 29053 31171 29056
rect 31113 29047 31171 29053
rect 3418 28976 3424 29028
rect 3476 29016 3482 29028
rect 25332 29016 25360 29047
rect 31754 29044 31760 29056
rect 31812 29044 31818 29096
rect 32214 29084 32220 29096
rect 32175 29056 32220 29084
rect 32214 29044 32220 29056
rect 32272 29044 32278 29096
rect 37366 29084 37372 29096
rect 37327 29056 37372 29084
rect 37366 29044 37372 29056
rect 37424 29044 37430 29096
rect 3476 28988 25360 29016
rect 3476 28976 3482 28988
rect 30834 28976 30840 29028
rect 30892 29016 30898 29028
rect 31021 29019 31079 29025
rect 31021 29016 31033 29019
rect 30892 28988 31033 29016
rect 30892 28976 30898 28988
rect 31021 28985 31033 28988
rect 31067 28985 31079 29019
rect 33502 29016 33508 29028
rect 33463 28988 33508 29016
rect 31021 28979 31079 28985
rect 33502 28976 33508 28988
rect 33560 28976 33566 29028
rect 36722 28976 36728 29028
rect 36780 29016 36786 29028
rect 36998 29016 37004 29028
rect 36780 28988 37004 29016
rect 36780 28976 36786 28988
rect 36998 28976 37004 28988
rect 37056 29016 37062 29028
rect 38580 29016 38608 29124
rect 38657 29121 38669 29124
rect 38703 29121 38715 29155
rect 38838 29152 38844 29164
rect 38799 29124 38844 29152
rect 38657 29115 38715 29121
rect 38838 29112 38844 29124
rect 38896 29112 38902 29164
rect 38933 29155 38991 29161
rect 38933 29121 38945 29155
rect 38979 29121 38991 29155
rect 39316 29150 39344 29260
rect 39592 29232 39620 29260
rect 42610 29248 42616 29260
rect 42668 29248 42674 29300
rect 43346 29288 43352 29300
rect 43307 29260 43352 29288
rect 43346 29248 43352 29260
rect 43404 29248 43410 29300
rect 43625 29291 43683 29297
rect 43625 29257 43637 29291
rect 43671 29288 43683 29291
rect 44266 29288 44272 29300
rect 43671 29260 44272 29288
rect 43671 29257 43683 29260
rect 43625 29251 43683 29257
rect 44266 29248 44272 29260
rect 44324 29248 44330 29300
rect 49970 29288 49976 29300
rect 49931 29260 49976 29288
rect 49970 29248 49976 29260
rect 50028 29248 50034 29300
rect 50614 29248 50620 29300
rect 50672 29288 50678 29300
rect 50801 29291 50859 29297
rect 50801 29288 50813 29291
rect 50672 29260 50813 29288
rect 50672 29248 50678 29260
rect 50801 29257 50813 29260
rect 50847 29257 50859 29291
rect 50801 29251 50859 29257
rect 50982 29248 50988 29300
rect 51040 29288 51046 29300
rect 51810 29288 51816 29300
rect 51040 29260 51085 29288
rect 51771 29260 51816 29288
rect 51040 29248 51046 29260
rect 51810 29248 51816 29260
rect 51868 29248 51874 29300
rect 52733 29291 52791 29297
rect 52733 29257 52745 29291
rect 52779 29288 52791 29291
rect 54386 29288 54392 29300
rect 52779 29260 54392 29288
rect 52779 29257 52791 29260
rect 52733 29251 52791 29257
rect 39574 29180 39580 29232
rect 39632 29220 39638 29232
rect 40773 29223 40831 29229
rect 40773 29220 40785 29223
rect 39632 29192 40785 29220
rect 39632 29180 39638 29192
rect 40773 29189 40785 29192
rect 40819 29189 40831 29223
rect 43257 29223 43315 29229
rect 43257 29220 43269 29223
rect 40773 29183 40831 29189
rect 42720 29192 43269 29220
rect 42720 29164 42748 29192
rect 43257 29189 43269 29192
rect 43303 29189 43315 29223
rect 43257 29183 43315 29189
rect 43438 29180 43444 29232
rect 43496 29220 43502 29232
rect 48682 29220 48688 29232
rect 43496 29192 48688 29220
rect 43496 29180 43502 29192
rect 48682 29180 48688 29192
rect 48740 29220 48746 29232
rect 49418 29220 49424 29232
rect 48740 29192 49424 29220
rect 48740 29180 48746 29192
rect 49418 29180 49424 29192
rect 49476 29220 49482 29232
rect 49476 29192 50752 29220
rect 49476 29180 49482 29192
rect 39393 29155 39451 29161
rect 39393 29150 39405 29155
rect 39316 29122 39405 29150
rect 38933 29115 38991 29121
rect 39393 29121 39405 29122
rect 39439 29121 39451 29155
rect 40586 29152 40592 29164
rect 39393 29115 39451 29121
rect 39592 29124 40592 29152
rect 38948 29084 38976 29115
rect 39592 29084 39620 29124
rect 40586 29112 40592 29124
rect 40644 29112 40650 29164
rect 40681 29155 40739 29161
rect 40681 29121 40693 29155
rect 40727 29152 40739 29155
rect 40954 29152 40960 29164
rect 40727 29124 40960 29152
rect 40727 29121 40739 29124
rect 40681 29115 40739 29121
rect 40954 29112 40960 29124
rect 41012 29112 41018 29164
rect 42426 29112 42432 29164
rect 42484 29152 42490 29164
rect 42521 29155 42579 29161
rect 42521 29152 42533 29155
rect 42484 29124 42533 29152
rect 42484 29112 42490 29124
rect 42521 29121 42533 29124
rect 42567 29121 42579 29155
rect 42702 29152 42708 29164
rect 42663 29124 42708 29152
rect 42521 29115 42579 29121
rect 38948 29056 39620 29084
rect 39669 29087 39727 29093
rect 39669 29053 39681 29087
rect 39715 29053 39727 29087
rect 42536 29084 42564 29115
rect 42702 29112 42708 29124
rect 42760 29112 42766 29164
rect 43162 29152 43168 29164
rect 43075 29124 43168 29152
rect 43162 29112 43168 29124
rect 43220 29152 43226 29164
rect 43625 29155 43683 29161
rect 43220 29124 43392 29152
rect 43220 29112 43226 29124
rect 43364 29084 43392 29124
rect 43625 29121 43637 29155
rect 43671 29152 43683 29155
rect 44174 29152 44180 29164
rect 43671 29124 44180 29152
rect 43671 29121 43683 29124
rect 43625 29115 43683 29121
rect 44174 29112 44180 29124
rect 44232 29112 44238 29164
rect 45925 29155 45983 29161
rect 45925 29121 45937 29155
rect 45971 29121 45983 29155
rect 45925 29115 45983 29121
rect 46109 29155 46167 29161
rect 46109 29121 46121 29155
rect 46155 29152 46167 29155
rect 46658 29152 46664 29164
rect 46155 29124 46664 29152
rect 46155 29121 46167 29124
rect 46109 29115 46167 29121
rect 42536 29056 43392 29084
rect 39669 29047 39727 29053
rect 37056 28988 38608 29016
rect 37056 28976 37062 28988
rect 38654 28976 38660 29028
rect 38712 29016 38718 29028
rect 39684 29016 39712 29047
rect 41138 29016 41144 29028
rect 38712 28988 41144 29016
rect 38712 28976 38718 28988
rect 41138 28976 41144 28988
rect 41196 28976 41202 29028
rect 43364 29016 43392 29056
rect 43487 29087 43545 29093
rect 43487 29053 43499 29087
rect 43533 29084 43545 29087
rect 43990 29084 43996 29096
rect 43533 29056 43996 29084
rect 43533 29053 43545 29056
rect 43487 29047 43545 29053
rect 43990 29044 43996 29056
rect 44048 29044 44054 29096
rect 45940 29084 45968 29115
rect 46658 29112 46664 29124
rect 46716 29152 46722 29164
rect 49786 29152 49792 29164
rect 46716 29124 49792 29152
rect 46716 29112 46722 29124
rect 49786 29112 49792 29124
rect 49844 29112 49850 29164
rect 49878 29112 49884 29164
rect 49936 29152 49942 29164
rect 50617 29155 50675 29161
rect 50617 29152 50629 29155
rect 49936 29124 50629 29152
rect 49936 29112 49942 29124
rect 50617 29121 50629 29124
rect 50663 29121 50675 29155
rect 50724 29152 50752 29192
rect 52454 29180 52460 29232
rect 52512 29220 52518 29232
rect 52512 29192 53144 29220
rect 52512 29180 52518 29192
rect 50893 29155 50951 29161
rect 50893 29152 50905 29155
rect 50724 29124 50905 29152
rect 50617 29115 50675 29121
rect 50893 29121 50905 29124
rect 50939 29121 50951 29155
rect 51442 29152 51448 29164
rect 50893 29115 50951 29121
rect 51108 29124 51448 29152
rect 46474 29084 46480 29096
rect 45940 29056 46480 29084
rect 46474 29044 46480 29056
rect 46532 29044 46538 29096
rect 50062 29044 50068 29096
rect 50120 29084 50126 29096
rect 50982 29084 50988 29096
rect 50120 29056 50988 29084
rect 50120 29044 50126 29056
rect 50982 29044 50988 29056
rect 51040 29044 51046 29096
rect 45646 29016 45652 29028
rect 43364 28988 45652 29016
rect 45646 28976 45652 28988
rect 45704 28976 45710 29028
rect 50614 28976 50620 29028
rect 50672 29016 50678 29028
rect 51108 29016 51136 29124
rect 51442 29112 51448 29124
rect 51500 29152 51506 29164
rect 53116 29161 53144 29192
rect 54128 29161 54156 29260
rect 54386 29248 54392 29260
rect 54444 29248 54450 29300
rect 54481 29291 54539 29297
rect 54481 29257 54493 29291
rect 54527 29288 54539 29291
rect 54754 29288 54760 29300
rect 54527 29260 54760 29288
rect 54527 29257 54539 29260
rect 54481 29251 54539 29257
rect 54754 29248 54760 29260
rect 54812 29248 54818 29300
rect 51721 29155 51779 29161
rect 51721 29152 51733 29155
rect 51500 29124 51733 29152
rect 51500 29112 51506 29124
rect 51721 29121 51733 29124
rect 51767 29121 51779 29155
rect 51721 29115 51779 29121
rect 53101 29155 53159 29161
rect 53101 29121 53113 29155
rect 53147 29121 53159 29155
rect 53101 29115 53159 29121
rect 54113 29155 54171 29161
rect 54113 29121 54125 29155
rect 54159 29121 54171 29155
rect 54113 29115 54171 29121
rect 52914 29084 52920 29096
rect 52875 29056 52920 29084
rect 52914 29044 52920 29056
rect 52972 29044 52978 29096
rect 53006 29044 53012 29096
rect 53064 29084 53070 29096
rect 53193 29087 53251 29093
rect 53064 29056 53109 29084
rect 53064 29044 53070 29056
rect 53193 29053 53205 29087
rect 53239 29053 53251 29087
rect 54018 29084 54024 29096
rect 53979 29056 54024 29084
rect 53193 29047 53251 29053
rect 50672 28988 51136 29016
rect 51169 29019 51227 29025
rect 50672 28976 50678 28988
rect 51169 28985 51181 29019
rect 51215 29016 51227 29019
rect 52822 29016 52828 29028
rect 51215 28988 52828 29016
rect 51215 28985 51227 28988
rect 51169 28979 51227 28985
rect 52822 28976 52828 28988
rect 52880 29016 52886 29028
rect 53208 29016 53236 29047
rect 54018 29044 54024 29056
rect 54076 29044 54082 29096
rect 52880 28988 53236 29016
rect 52880 28976 52886 28988
rect 30653 28951 30711 28957
rect 30653 28917 30665 28951
rect 30699 28948 30711 28951
rect 31478 28948 31484 28960
rect 30699 28920 31484 28948
rect 30699 28917 30711 28920
rect 30653 28911 30711 28917
rect 31478 28908 31484 28920
rect 31536 28908 31542 28960
rect 32306 28948 32312 28960
rect 32267 28920 32312 28948
rect 32306 28908 32312 28920
rect 32364 28908 32370 28960
rect 37458 28948 37464 28960
rect 37419 28920 37464 28948
rect 37458 28908 37464 28920
rect 37516 28908 37522 28960
rect 37645 28951 37703 28957
rect 37645 28917 37657 28951
rect 37691 28948 37703 28951
rect 38010 28948 38016 28960
rect 37691 28920 38016 28948
rect 37691 28917 37703 28920
rect 37645 28911 37703 28917
rect 38010 28908 38016 28920
rect 38068 28908 38074 28960
rect 38286 28948 38292 28960
rect 38247 28920 38292 28948
rect 38286 28908 38292 28920
rect 38344 28908 38350 28960
rect 40862 28908 40868 28960
rect 40920 28948 40926 28960
rect 42518 28948 42524 28960
rect 40920 28920 42524 28948
rect 40920 28908 40926 28920
rect 42518 28908 42524 28920
rect 42576 28908 42582 28960
rect 45922 28948 45928 28960
rect 45883 28920 45928 28948
rect 45922 28908 45928 28920
rect 45980 28908 45986 28960
rect 46014 28908 46020 28960
rect 46072 28948 46078 28960
rect 48498 28948 48504 28960
rect 46072 28920 48504 28948
rect 46072 28908 46078 28920
rect 48498 28908 48504 28920
rect 48556 28908 48562 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 25222 28744 25228 28756
rect 25183 28716 25228 28744
rect 25222 28704 25228 28716
rect 25280 28704 25286 28756
rect 27157 28747 27215 28753
rect 27157 28713 27169 28747
rect 27203 28744 27215 28747
rect 27246 28744 27252 28756
rect 27203 28716 27252 28744
rect 27203 28713 27215 28716
rect 27157 28707 27215 28713
rect 27246 28704 27252 28716
rect 27304 28704 27310 28756
rect 28258 28704 28264 28756
rect 28316 28744 28322 28756
rect 40862 28744 40868 28756
rect 28316 28716 40868 28744
rect 28316 28704 28322 28716
rect 40862 28704 40868 28716
rect 40920 28704 40926 28756
rect 47486 28744 47492 28756
rect 42444 28716 47492 28744
rect 28813 28679 28871 28685
rect 28813 28676 28825 28679
rect 28736 28648 28825 28676
rect 28534 28608 28540 28620
rect 28495 28580 28540 28608
rect 28534 28568 28540 28580
rect 28592 28568 28598 28620
rect 25133 28543 25191 28549
rect 25133 28509 25145 28543
rect 25179 28509 25191 28543
rect 25133 28503 25191 28509
rect 24854 28364 24860 28416
rect 24912 28404 24918 28416
rect 25148 28404 25176 28503
rect 26142 28500 26148 28552
rect 26200 28540 26206 28552
rect 27154 28540 27160 28552
rect 26200 28512 27160 28540
rect 26200 28500 26206 28512
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 27338 28540 27344 28552
rect 27299 28512 27344 28540
rect 27338 28500 27344 28512
rect 27396 28500 27402 28552
rect 28552 28472 28580 28568
rect 28736 28540 28764 28648
rect 28813 28645 28825 28648
rect 28859 28645 28871 28679
rect 28813 28639 28871 28645
rect 28997 28679 29055 28685
rect 28997 28645 29009 28679
rect 29043 28676 29055 28679
rect 32306 28676 32312 28688
rect 29043 28648 32312 28676
rect 29043 28645 29055 28648
rect 28997 28639 29055 28645
rect 32306 28636 32312 28648
rect 32364 28676 32370 28688
rect 32364 28648 33456 28676
rect 32364 28636 32370 28648
rect 29549 28611 29607 28617
rect 29549 28577 29561 28611
rect 29595 28577 29607 28611
rect 29549 28571 29607 28577
rect 31297 28611 31355 28617
rect 31297 28577 31309 28611
rect 31343 28608 31355 28611
rect 31938 28608 31944 28620
rect 31343 28580 31944 28608
rect 31343 28577 31355 28580
rect 31297 28571 31355 28577
rect 28994 28540 29000 28552
rect 28736 28512 29000 28540
rect 28994 28500 29000 28512
rect 29052 28500 29058 28552
rect 29564 28472 29592 28571
rect 31938 28568 31944 28580
rect 31996 28608 32002 28620
rect 31996 28580 33088 28608
rect 31996 28568 32002 28580
rect 29822 28540 29828 28552
rect 29783 28512 29828 28540
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 31110 28500 31116 28552
rect 31168 28540 31174 28552
rect 31573 28543 31631 28549
rect 31573 28540 31585 28543
rect 31168 28512 31585 28540
rect 31168 28500 31174 28512
rect 31573 28509 31585 28512
rect 31619 28509 31631 28543
rect 32674 28540 32680 28552
rect 32635 28512 32680 28540
rect 31573 28503 31631 28509
rect 32674 28500 32680 28512
rect 32732 28500 32738 28552
rect 32858 28540 32864 28552
rect 32819 28512 32864 28540
rect 32858 28500 32864 28512
rect 32916 28500 32922 28552
rect 28552 28444 29592 28472
rect 30374 28432 30380 28484
rect 30432 28472 30438 28484
rect 32953 28475 33011 28481
rect 32953 28472 32965 28475
rect 30432 28444 32965 28472
rect 30432 28432 30438 28444
rect 32953 28441 32965 28444
rect 32999 28441 33011 28475
rect 33060 28472 33088 28580
rect 33428 28549 33456 28648
rect 36814 28636 36820 28688
rect 36872 28676 36878 28688
rect 36909 28679 36967 28685
rect 36909 28676 36921 28679
rect 36872 28648 36921 28676
rect 36872 28636 36878 28648
rect 36909 28645 36921 28648
rect 36955 28645 36967 28679
rect 40770 28676 40776 28688
rect 36909 28639 36967 28645
rect 37476 28648 40776 28676
rect 34698 28608 34704 28620
rect 34659 28580 34704 28608
rect 34698 28568 34704 28580
rect 34756 28568 34762 28620
rect 35802 28568 35808 28620
rect 35860 28608 35866 28620
rect 37476 28608 37504 28648
rect 40770 28636 40776 28648
rect 40828 28636 40834 28688
rect 41325 28679 41383 28685
rect 41325 28645 41337 28679
rect 41371 28645 41383 28679
rect 41325 28639 41383 28645
rect 35860 28580 37504 28608
rect 37553 28611 37611 28617
rect 35860 28568 35866 28580
rect 37553 28577 37565 28611
rect 37599 28608 37611 28611
rect 41340 28608 41368 28639
rect 42444 28608 42472 28716
rect 47486 28704 47492 28716
rect 47544 28704 47550 28756
rect 47946 28704 47952 28756
rect 48004 28744 48010 28756
rect 48409 28747 48467 28753
rect 48409 28744 48421 28747
rect 48004 28716 48421 28744
rect 48004 28704 48010 28716
rect 48409 28713 48421 28716
rect 48455 28713 48467 28747
rect 48774 28744 48780 28756
rect 48735 28716 48780 28744
rect 48409 28707 48467 28713
rect 48774 28704 48780 28716
rect 48832 28704 48838 28756
rect 52822 28744 52828 28756
rect 52783 28716 52828 28744
rect 52822 28704 52828 28716
rect 52880 28704 52886 28756
rect 53006 28704 53012 28756
rect 53064 28744 53070 28756
rect 53561 28747 53619 28753
rect 53561 28744 53573 28747
rect 53064 28716 53573 28744
rect 53064 28704 53070 28716
rect 53561 28713 53573 28716
rect 53607 28713 53619 28747
rect 53561 28707 53619 28713
rect 54665 28747 54723 28753
rect 54665 28713 54677 28747
rect 54711 28744 54723 28747
rect 55306 28744 55312 28756
rect 54711 28716 55312 28744
rect 54711 28713 54723 28716
rect 54665 28707 54723 28713
rect 55306 28704 55312 28716
rect 55364 28704 55370 28756
rect 42518 28636 42524 28688
rect 42576 28676 42582 28688
rect 55214 28676 55220 28688
rect 42576 28648 55220 28676
rect 42576 28636 42582 28648
rect 55214 28636 55220 28648
rect 55272 28636 55278 28688
rect 37599 28580 41276 28608
rect 41340 28580 42472 28608
rect 37599 28577 37611 28580
rect 37553 28571 37611 28577
rect 33413 28543 33471 28549
rect 33413 28509 33425 28543
rect 33459 28509 33471 28543
rect 33413 28503 33471 28509
rect 33597 28543 33655 28549
rect 33597 28509 33609 28543
rect 33643 28509 33655 28543
rect 37734 28540 37740 28552
rect 37695 28512 37740 28540
rect 33597 28503 33655 28509
rect 33612 28472 33640 28503
rect 37734 28500 37740 28512
rect 37792 28500 37798 28552
rect 38010 28540 38016 28552
rect 37971 28512 38016 28540
rect 38010 28500 38016 28512
rect 38068 28500 38074 28552
rect 38841 28543 38899 28549
rect 38841 28509 38853 28543
rect 38887 28540 38899 28543
rect 38930 28540 38936 28552
rect 38887 28512 38936 28540
rect 38887 28509 38899 28512
rect 38841 28503 38899 28509
rect 38930 28500 38936 28512
rect 38988 28500 38994 28552
rect 39025 28543 39083 28549
rect 39025 28509 39037 28543
rect 39071 28540 39083 28543
rect 40954 28540 40960 28552
rect 39071 28512 40960 28540
rect 39071 28509 39083 28512
rect 39025 28503 39083 28509
rect 33060 28444 33640 28472
rect 34968 28475 35026 28481
rect 32953 28435 33011 28441
rect 34968 28441 34980 28475
rect 35014 28472 35026 28475
rect 35618 28472 35624 28484
rect 35014 28444 35624 28472
rect 35014 28441 35026 28444
rect 34968 28435 35026 28441
rect 35618 28432 35624 28444
rect 35676 28432 35682 28484
rect 36725 28475 36783 28481
rect 36725 28441 36737 28475
rect 36771 28472 36783 28475
rect 37182 28472 37188 28484
rect 36771 28444 37188 28472
rect 36771 28441 36783 28444
rect 36725 28435 36783 28441
rect 37182 28432 37188 28444
rect 37240 28432 37246 28484
rect 37274 28432 37280 28484
rect 37332 28472 37338 28484
rect 39040 28472 39068 28503
rect 40954 28500 40960 28512
rect 41012 28500 41018 28552
rect 41138 28540 41144 28552
rect 41099 28512 41144 28540
rect 41138 28500 41144 28512
rect 41196 28500 41202 28552
rect 41248 28540 41276 28580
rect 42886 28568 42892 28620
rect 42944 28608 42950 28620
rect 43346 28608 43352 28620
rect 42944 28580 43352 28608
rect 42944 28568 42950 28580
rect 43346 28568 43352 28580
rect 43404 28608 43410 28620
rect 45830 28608 45836 28620
rect 43404 28580 43944 28608
rect 43404 28568 43410 28580
rect 41782 28540 41788 28552
rect 41248 28512 41788 28540
rect 41782 28500 41788 28512
rect 41840 28500 41846 28552
rect 43714 28540 43720 28552
rect 43675 28512 43720 28540
rect 43714 28500 43720 28512
rect 43772 28500 43778 28552
rect 43916 28549 43944 28580
rect 45168 28580 45836 28608
rect 43901 28543 43959 28549
rect 43901 28509 43913 28543
rect 43947 28509 43959 28543
rect 45002 28540 45008 28552
rect 44963 28512 45008 28540
rect 43901 28503 43959 28509
rect 45002 28500 45008 28512
rect 45060 28500 45066 28552
rect 45168 28549 45196 28580
rect 45830 28568 45836 28580
rect 45888 28568 45894 28620
rect 47946 28608 47952 28620
rect 46676 28580 47952 28608
rect 45554 28549 45560 28552
rect 45153 28543 45211 28549
rect 45153 28509 45165 28543
rect 45199 28509 45211 28543
rect 45153 28503 45211 28509
rect 45509 28543 45560 28549
rect 45509 28509 45521 28543
rect 45555 28509 45560 28543
rect 45509 28503 45560 28509
rect 45554 28500 45560 28503
rect 45612 28500 45618 28552
rect 46676 28549 46704 28580
rect 47946 28568 47952 28580
rect 48004 28568 48010 28620
rect 51813 28611 51871 28617
rect 51813 28577 51825 28611
rect 51859 28608 51871 28611
rect 57790 28608 57796 28620
rect 51859 28580 54524 28608
rect 57751 28580 57796 28608
rect 51859 28577 51871 28580
rect 51813 28571 51871 28577
rect 46661 28543 46719 28549
rect 46661 28509 46673 28543
rect 46707 28509 46719 28543
rect 46661 28503 46719 28509
rect 46937 28543 46995 28549
rect 46937 28509 46949 28543
rect 46983 28509 46995 28543
rect 46937 28503 46995 28509
rect 37332 28444 39068 28472
rect 37332 28432 37338 28444
rect 40218 28432 40224 28484
rect 40276 28472 40282 28484
rect 40313 28475 40371 28481
rect 40313 28472 40325 28475
rect 40276 28444 40325 28472
rect 40276 28432 40282 28444
rect 40313 28441 40325 28444
rect 40359 28441 40371 28475
rect 40678 28472 40684 28484
rect 40639 28444 40684 28472
rect 40313 28435 40371 28441
rect 40678 28432 40684 28444
rect 40736 28432 40742 28484
rect 40770 28432 40776 28484
rect 40828 28472 40834 28484
rect 45278 28472 45284 28484
rect 40828 28444 44220 28472
rect 45239 28444 45284 28472
rect 40828 28432 40834 28444
rect 33134 28404 33140 28416
rect 24912 28376 33140 28404
rect 24912 28364 24918 28376
rect 33134 28364 33140 28376
rect 33192 28364 33198 28416
rect 33502 28404 33508 28416
rect 33463 28376 33508 28404
rect 33502 28364 33508 28376
rect 33560 28364 33566 28416
rect 36081 28407 36139 28413
rect 36081 28373 36093 28407
rect 36127 28404 36139 28407
rect 36170 28404 36176 28416
rect 36127 28376 36176 28404
rect 36127 28373 36139 28376
rect 36081 28367 36139 28373
rect 36170 28364 36176 28376
rect 36228 28364 36234 28416
rect 37921 28407 37979 28413
rect 37921 28373 37933 28407
rect 37967 28404 37979 28407
rect 38102 28404 38108 28416
rect 37967 28376 38108 28404
rect 37967 28373 37979 28376
rect 37921 28367 37979 28373
rect 38102 28364 38108 28376
rect 38160 28364 38166 28416
rect 43898 28404 43904 28416
rect 43859 28376 43904 28404
rect 43898 28364 43904 28376
rect 43956 28364 43962 28416
rect 44192 28404 44220 28444
rect 45278 28432 45284 28444
rect 45336 28432 45342 28484
rect 45370 28432 45376 28484
rect 45428 28481 45434 28484
rect 45428 28472 45439 28481
rect 46014 28472 46020 28484
rect 45428 28444 46020 28472
rect 45428 28435 45439 28444
rect 45428 28432 45434 28435
rect 46014 28432 46020 28444
rect 46072 28432 46078 28484
rect 46952 28472 46980 28503
rect 47210 28500 47216 28552
rect 47268 28540 47274 28552
rect 47581 28543 47639 28549
rect 47581 28540 47593 28543
rect 47268 28512 47593 28540
rect 47268 28500 47274 28512
rect 47581 28509 47593 28512
rect 47627 28509 47639 28543
rect 47762 28540 47768 28552
rect 47723 28512 47768 28540
rect 47581 28503 47639 28509
rect 47762 28500 47768 28512
rect 47820 28500 47826 28552
rect 47854 28500 47860 28552
rect 47912 28540 47918 28552
rect 48317 28543 48375 28549
rect 47912 28512 47957 28540
rect 47912 28500 47918 28512
rect 48317 28509 48329 28543
rect 48363 28509 48375 28543
rect 50154 28540 50160 28552
rect 50115 28512 50160 28540
rect 48317 28503 48375 28509
rect 47397 28475 47455 28481
rect 47397 28472 47409 28475
rect 46952 28444 47409 28472
rect 47397 28441 47409 28444
rect 47443 28472 47455 28475
rect 48332 28472 48360 28503
rect 50154 28500 50160 28512
rect 50212 28500 50218 28552
rect 50433 28543 50491 28549
rect 50433 28509 50445 28543
rect 50479 28540 50491 28543
rect 50614 28540 50620 28552
rect 50479 28512 50620 28540
rect 50479 28509 50491 28512
rect 50433 28503 50491 28509
rect 50614 28500 50620 28512
rect 50672 28500 50678 28552
rect 51445 28543 51503 28549
rect 51445 28509 51457 28543
rect 51491 28540 51503 28543
rect 51902 28540 51908 28552
rect 51491 28512 51908 28540
rect 51491 28509 51503 28512
rect 51445 28503 51503 28509
rect 51902 28500 51908 28512
rect 51960 28500 51966 28552
rect 52454 28540 52460 28552
rect 52415 28512 52460 28540
rect 52454 28500 52460 28512
rect 52512 28500 52518 28552
rect 52914 28500 52920 28552
rect 52972 28540 52978 28552
rect 54496 28549 54524 28580
rect 57790 28568 57796 28580
rect 57848 28568 57854 28620
rect 54481 28543 54539 28549
rect 52972 28512 53017 28540
rect 52972 28500 52978 28512
rect 54481 28509 54493 28543
rect 54527 28540 54539 28543
rect 54662 28540 54668 28552
rect 54527 28512 54668 28540
rect 54527 28509 54539 28512
rect 54481 28503 54539 28509
rect 54662 28500 54668 28512
rect 54720 28500 54726 28552
rect 56318 28540 56324 28552
rect 56279 28512 56324 28540
rect 56318 28500 56324 28512
rect 56376 28500 56382 28552
rect 51626 28472 51632 28484
rect 47443 28444 48360 28472
rect 51587 28444 51632 28472
rect 47443 28441 47455 28444
rect 47397 28435 47455 28441
rect 51626 28432 51632 28444
rect 51684 28432 51690 28484
rect 53190 28472 53196 28484
rect 52288 28444 53196 28472
rect 45186 28404 45192 28416
rect 44192 28376 45192 28404
rect 45186 28364 45192 28376
rect 45244 28364 45250 28416
rect 45646 28364 45652 28416
rect 45704 28404 45710 28416
rect 45704 28376 45749 28404
rect 45704 28364 45710 28376
rect 45830 28364 45836 28416
rect 45888 28404 45894 28416
rect 46477 28407 46535 28413
rect 46477 28404 46489 28407
rect 45888 28376 46489 28404
rect 45888 28364 45894 28376
rect 46477 28373 46489 28376
rect 46523 28373 46535 28407
rect 46477 28367 46535 28373
rect 46845 28407 46903 28413
rect 46845 28373 46857 28407
rect 46891 28404 46903 28407
rect 47578 28404 47584 28416
rect 46891 28376 47584 28404
rect 46891 28373 46903 28376
rect 46845 28367 46903 28373
rect 47578 28364 47584 28376
rect 47636 28364 47642 28416
rect 52288 28413 52316 28444
rect 53190 28432 53196 28444
rect 53248 28432 53254 28484
rect 53469 28475 53527 28481
rect 53469 28441 53481 28475
rect 53515 28441 53527 28475
rect 53469 28435 53527 28441
rect 54297 28475 54355 28481
rect 54297 28441 54309 28475
rect 54343 28472 54355 28475
rect 54386 28472 54392 28484
rect 54343 28444 54392 28472
rect 54343 28441 54355 28444
rect 54297 28435 54355 28441
rect 52273 28407 52331 28413
rect 52273 28373 52285 28407
rect 52319 28373 52331 28407
rect 52273 28367 52331 28373
rect 52362 28364 52368 28416
rect 52420 28404 52426 28416
rect 52457 28407 52515 28413
rect 52457 28404 52469 28407
rect 52420 28376 52469 28404
rect 52420 28364 52426 28376
rect 52457 28373 52469 28376
rect 52503 28404 52515 28407
rect 53484 28404 53512 28435
rect 54386 28432 54392 28444
rect 54444 28432 54450 28484
rect 56505 28475 56563 28481
rect 56505 28441 56517 28475
rect 56551 28472 56563 28475
rect 56962 28472 56968 28484
rect 56551 28444 56968 28472
rect 56551 28441 56563 28444
rect 56505 28435 56563 28441
rect 56962 28432 56968 28444
rect 57020 28432 57026 28484
rect 52503 28376 53512 28404
rect 52503 28373 52515 28376
rect 52457 28367 52515 28373
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 29003 28203 29061 28209
rect 29003 28169 29015 28203
rect 29049 28200 29061 28203
rect 31018 28200 31024 28212
rect 29049 28172 31024 28200
rect 29049 28169 29061 28172
rect 29003 28163 29061 28169
rect 31018 28160 31024 28172
rect 31076 28160 31082 28212
rect 31570 28160 31576 28212
rect 31628 28200 31634 28212
rect 31628 28172 32628 28200
rect 31628 28160 31634 28172
rect 29089 28135 29147 28141
rect 29089 28101 29101 28135
rect 29135 28132 29147 28135
rect 30929 28135 30987 28141
rect 29135 28104 29592 28132
rect 29135 28101 29147 28104
rect 29089 28095 29147 28101
rect 28810 28024 28816 28076
rect 28868 28064 28874 28076
rect 28905 28067 28963 28073
rect 28905 28064 28917 28067
rect 28868 28036 28917 28064
rect 28868 28024 28874 28036
rect 28905 28033 28917 28036
rect 28951 28033 28963 28067
rect 28905 28027 28963 28033
rect 29181 28067 29239 28073
rect 29181 28033 29193 28067
rect 29227 28064 29239 28067
rect 29270 28064 29276 28076
rect 29227 28036 29276 28064
rect 29227 28033 29239 28036
rect 29181 28027 29239 28033
rect 29270 28024 29276 28036
rect 29328 28024 29334 28076
rect 29564 28064 29592 28104
rect 30929 28101 30941 28135
rect 30975 28132 30987 28135
rect 32600 28132 32628 28172
rect 32674 28160 32680 28212
rect 32732 28200 32738 28212
rect 33321 28203 33379 28209
rect 33321 28200 33333 28203
rect 32732 28172 33333 28200
rect 32732 28160 32738 28172
rect 33321 28169 33333 28172
rect 33367 28169 33379 28203
rect 33321 28163 33379 28169
rect 36449 28203 36507 28209
rect 36449 28169 36461 28203
rect 36495 28200 36507 28203
rect 38286 28200 38292 28212
rect 36495 28172 38292 28200
rect 36495 28169 36507 28172
rect 36449 28163 36507 28169
rect 38286 28160 38292 28172
rect 38344 28160 38350 28212
rect 39206 28160 39212 28212
rect 39264 28160 39270 28212
rect 43346 28200 43352 28212
rect 43307 28172 43352 28200
rect 43346 28160 43352 28172
rect 43404 28160 43410 28212
rect 44358 28200 44364 28212
rect 44319 28172 44364 28200
rect 44358 28160 44364 28172
rect 44416 28160 44422 28212
rect 44913 28203 44971 28209
rect 44913 28169 44925 28203
rect 44959 28200 44971 28203
rect 45094 28200 45100 28212
rect 44959 28172 45100 28200
rect 44959 28169 44971 28172
rect 44913 28163 44971 28169
rect 45094 28160 45100 28172
rect 45152 28200 45158 28212
rect 45554 28200 45560 28212
rect 45152 28172 45560 28200
rect 45152 28160 45158 28172
rect 45554 28160 45560 28172
rect 45612 28160 45618 28212
rect 46017 28203 46075 28209
rect 46017 28169 46029 28203
rect 46063 28200 46075 28203
rect 46106 28200 46112 28212
rect 46063 28172 46112 28200
rect 46063 28169 46075 28172
rect 46017 28163 46075 28169
rect 46106 28160 46112 28172
rect 46164 28160 46170 28212
rect 47946 28200 47952 28212
rect 47907 28172 47952 28200
rect 47946 28160 47952 28172
rect 48004 28160 48010 28212
rect 48314 28160 48320 28212
rect 48372 28200 48378 28212
rect 49602 28200 49608 28212
rect 48372 28172 49608 28200
rect 48372 28160 48378 28172
rect 49602 28160 49608 28172
rect 49660 28160 49666 28212
rect 50062 28160 50068 28212
rect 50120 28200 50126 28212
rect 50295 28203 50353 28209
rect 50295 28200 50307 28203
rect 50120 28172 50307 28200
rect 50120 28160 50126 28172
rect 50295 28169 50307 28172
rect 50341 28169 50353 28203
rect 50295 28163 50353 28169
rect 53006 28160 53012 28212
rect 53064 28200 53070 28212
rect 53064 28172 53236 28200
rect 53064 28160 53070 28172
rect 33502 28132 33508 28144
rect 30975 28104 32174 28132
rect 32600 28104 33508 28132
rect 30975 28101 30987 28104
rect 30929 28095 30987 28101
rect 31202 28064 31208 28076
rect 29564 28036 31064 28064
rect 31163 28036 31208 28064
rect 28994 27956 29000 28008
rect 29052 27996 29058 28008
rect 29638 27996 29644 28008
rect 29052 27968 29644 27996
rect 29052 27956 29058 27968
rect 29638 27956 29644 27968
rect 29696 27956 29702 28008
rect 31036 27996 31064 28036
rect 31202 28024 31208 28036
rect 31260 28024 31266 28076
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28033 31355 28067
rect 31297 28027 31355 28033
rect 31389 28067 31447 28073
rect 31389 28033 31401 28067
rect 31435 28064 31447 28067
rect 31478 28064 31484 28076
rect 31435 28036 31484 28064
rect 31435 28033 31447 28036
rect 31389 28027 31447 28033
rect 31110 27996 31116 28008
rect 31023 27968 31116 27996
rect 31110 27956 31116 27968
rect 31168 27996 31174 28008
rect 31312 27996 31340 28027
rect 31478 28024 31484 28036
rect 31536 28024 31542 28076
rect 31570 28024 31576 28076
rect 31628 28064 31634 28076
rect 32146 28073 32174 28104
rect 32125 28067 32183 28073
rect 31628 28036 31673 28064
rect 31628 28024 31634 28036
rect 32125 28033 32137 28067
rect 32171 28033 32183 28067
rect 33042 28064 33048 28076
rect 33003 28036 33048 28064
rect 32125 28027 32183 28033
rect 33042 28024 33048 28036
rect 33100 28024 33106 28076
rect 32214 27996 32220 28008
rect 31168 27968 31340 27996
rect 32127 27968 32220 27996
rect 31168 27956 31174 27968
rect 32214 27956 32220 27968
rect 32272 27996 32278 28008
rect 32674 27996 32680 28008
rect 32272 27968 32680 27996
rect 32272 27956 32278 27968
rect 32674 27956 32680 27968
rect 32732 27956 32738 28008
rect 33336 28005 33364 28104
rect 33502 28092 33508 28104
rect 33560 28092 33566 28144
rect 34054 28141 34060 28144
rect 34048 28132 34060 28141
rect 34015 28104 34060 28132
rect 34048 28095 34060 28104
rect 34054 28092 34060 28095
rect 34112 28092 34118 28144
rect 36556 28104 37320 28132
rect 33778 28064 33784 28076
rect 33739 28036 33784 28064
rect 33778 28024 33784 28036
rect 33836 28024 33842 28076
rect 35713 28067 35771 28073
rect 35713 28033 35725 28067
rect 35759 28064 35771 28067
rect 36170 28064 36176 28076
rect 35759 28036 36176 28064
rect 35759 28033 35771 28036
rect 35713 28027 35771 28033
rect 36170 28024 36176 28036
rect 36228 28024 36234 28076
rect 36354 28064 36360 28076
rect 36315 28036 36360 28064
rect 36354 28024 36360 28036
rect 36412 28024 36418 28076
rect 36556 28005 36584 28104
rect 37292 28076 37320 28104
rect 37734 28092 37740 28144
rect 37792 28132 37798 28144
rect 39224 28132 39252 28160
rect 37792 28104 38608 28132
rect 39224 28104 39436 28132
rect 37792 28092 37798 28104
rect 36725 28067 36783 28073
rect 36725 28033 36737 28067
rect 36771 28033 36783 28067
rect 37274 28064 37280 28076
rect 37235 28036 37280 28064
rect 36725 28027 36783 28033
rect 33321 27999 33379 28005
rect 33321 27965 33333 27999
rect 33367 27965 33379 27999
rect 33321 27959 33379 27965
rect 36541 27999 36599 28005
rect 36541 27965 36553 27999
rect 36587 27965 36599 27999
rect 36740 27996 36768 28027
rect 37274 28024 37280 28036
rect 37332 28024 37338 28076
rect 37458 28024 37464 28076
rect 37516 28064 37522 28076
rect 37829 28067 37887 28073
rect 37829 28064 37841 28067
rect 37516 28036 37841 28064
rect 37516 28024 37522 28036
rect 37829 28033 37841 28036
rect 37875 28033 37887 28067
rect 37829 28027 37887 28033
rect 37844 27996 37872 28027
rect 37918 28024 37924 28076
rect 37976 28064 37982 28076
rect 38013 28067 38071 28073
rect 38013 28064 38025 28067
rect 37976 28036 38025 28064
rect 37976 28024 37982 28036
rect 38013 28033 38025 28036
rect 38059 28033 38071 28067
rect 38013 28027 38071 28033
rect 38378 28024 38384 28076
rect 38436 28064 38442 28076
rect 38580 28073 38608 28104
rect 38473 28067 38531 28073
rect 38473 28064 38485 28067
rect 38436 28036 38485 28064
rect 38436 28024 38442 28036
rect 38473 28033 38485 28036
rect 38519 28033 38531 28067
rect 38473 28027 38531 28033
rect 38565 28067 38623 28073
rect 38565 28033 38577 28067
rect 38611 28033 38623 28067
rect 39206 28064 39212 28076
rect 39167 28036 39212 28064
rect 38565 28027 38623 28033
rect 39206 28024 39212 28036
rect 39264 28024 39270 28076
rect 39408 28073 39436 28104
rect 40954 28092 40960 28144
rect 41012 28132 41018 28144
rect 41049 28135 41107 28141
rect 41049 28132 41061 28135
rect 41012 28104 41061 28132
rect 41012 28092 41018 28104
rect 41049 28101 41061 28104
rect 41095 28101 41107 28135
rect 41049 28095 41107 28101
rect 43438 28092 43444 28144
rect 43496 28132 43502 28144
rect 45370 28132 45376 28144
rect 43496 28104 45376 28132
rect 43496 28092 43502 28104
rect 45370 28092 45376 28104
rect 45428 28092 45434 28144
rect 47210 28092 47216 28144
rect 47268 28132 47274 28144
rect 47581 28135 47639 28141
rect 47581 28132 47593 28135
rect 47268 28104 47593 28132
rect 47268 28092 47274 28104
rect 47581 28101 47593 28104
rect 47627 28101 47639 28135
rect 47854 28132 47860 28144
rect 47581 28095 47639 28101
rect 47796 28101 47860 28132
rect 39393 28067 39451 28073
rect 39393 28033 39405 28067
rect 39439 28033 39451 28067
rect 39393 28027 39451 28033
rect 43165 28067 43223 28073
rect 43165 28033 43177 28067
rect 43211 28033 43223 28067
rect 43165 28027 43223 28033
rect 39301 27999 39359 28005
rect 39301 27996 39313 27999
rect 36740 27968 37780 27996
rect 37844 27968 39313 27996
rect 36541 27959 36599 27965
rect 29362 27888 29368 27940
rect 29420 27928 29426 27940
rect 29822 27928 29828 27940
rect 29420 27900 29828 27928
rect 29420 27888 29426 27900
rect 29822 27888 29828 27900
rect 29880 27928 29886 27940
rect 29917 27931 29975 27937
rect 29917 27928 29929 27931
rect 29880 27900 29929 27928
rect 29880 27888 29886 27900
rect 29917 27897 29929 27900
rect 29963 27897 29975 27931
rect 29917 27891 29975 27897
rect 30101 27931 30159 27937
rect 30101 27897 30113 27931
rect 30147 27928 30159 27931
rect 33137 27931 33195 27937
rect 33137 27928 33149 27931
rect 30147 27900 33149 27928
rect 30147 27897 30159 27900
rect 30101 27891 30159 27897
rect 33137 27897 33149 27900
rect 33183 27897 33195 27931
rect 33137 27891 33195 27897
rect 35805 27931 35863 27937
rect 35805 27897 35817 27931
rect 35851 27928 35863 27931
rect 37182 27928 37188 27940
rect 35851 27900 37188 27928
rect 35851 27897 35863 27900
rect 35805 27891 35863 27897
rect 28994 27820 29000 27872
rect 29052 27860 29058 27872
rect 29270 27860 29276 27872
rect 29052 27832 29276 27860
rect 29052 27820 29058 27832
rect 29270 27820 29276 27832
rect 29328 27860 29334 27872
rect 30116 27860 30144 27891
rect 37182 27888 37188 27900
rect 37240 27888 37246 27940
rect 37752 27928 37780 27968
rect 39301 27965 39313 27968
rect 39347 27965 39359 27999
rect 39301 27959 39359 27965
rect 39022 27928 39028 27940
rect 37752 27900 39028 27928
rect 39022 27888 39028 27900
rect 39080 27888 39086 27940
rect 32122 27860 32128 27872
rect 29328 27832 30144 27860
rect 32083 27832 32128 27860
rect 29328 27820 29334 27832
rect 32122 27820 32128 27832
rect 32180 27820 32186 27872
rect 32493 27863 32551 27869
rect 32493 27829 32505 27863
rect 32539 27860 32551 27863
rect 34422 27860 34428 27872
rect 32539 27832 34428 27860
rect 32539 27829 32551 27832
rect 32493 27823 32551 27829
rect 34422 27820 34428 27832
rect 34480 27820 34486 27872
rect 35161 27863 35219 27869
rect 35161 27829 35173 27863
rect 35207 27860 35219 27863
rect 36538 27860 36544 27872
rect 35207 27832 36544 27860
rect 35207 27829 35219 27832
rect 35161 27823 35219 27829
rect 36538 27820 36544 27832
rect 36596 27820 36602 27872
rect 36725 27863 36783 27869
rect 36725 27829 36737 27863
rect 36771 27860 36783 27863
rect 37734 27860 37740 27872
rect 36771 27832 37740 27860
rect 36771 27829 36783 27832
rect 36725 27823 36783 27829
rect 37734 27820 37740 27832
rect 37792 27820 37798 27872
rect 37826 27820 37832 27872
rect 37884 27860 37890 27872
rect 39408 27860 39436 28027
rect 43180 27928 43208 28027
rect 43254 28024 43260 28076
rect 43312 28064 43318 28076
rect 43349 28067 43407 28073
rect 43349 28064 43361 28067
rect 43312 28036 43361 28064
rect 43312 28024 43318 28036
rect 43349 28033 43361 28036
rect 43395 28033 43407 28067
rect 43349 28027 43407 28033
rect 43993 28067 44051 28073
rect 43993 28033 44005 28067
rect 44039 28064 44051 28067
rect 44726 28064 44732 28076
rect 44039 28036 44732 28064
rect 44039 28033 44051 28036
rect 43993 28027 44051 28033
rect 44726 28024 44732 28036
rect 44784 28024 44790 28076
rect 44821 28067 44879 28073
rect 44821 28033 44833 28067
rect 44867 28033 44879 28067
rect 44821 28027 44879 28033
rect 45649 28067 45707 28073
rect 45649 28033 45661 28067
rect 45695 28064 45707 28067
rect 46382 28064 46388 28076
rect 45695 28036 46388 28064
rect 45695 28033 45707 28036
rect 45649 28027 45707 28033
rect 43898 27996 43904 28008
rect 43859 27968 43904 27996
rect 43898 27956 43904 27968
rect 43956 27956 43962 28008
rect 44836 27928 44864 28027
rect 46382 28024 46388 28036
rect 46440 28024 46446 28076
rect 46474 28024 46480 28076
rect 46532 28064 46538 28076
rect 46532 28036 46577 28064
rect 46532 28024 46538 28036
rect 46658 28024 46664 28076
rect 46716 28064 46722 28076
rect 47796 28070 47823 28101
rect 47811 28067 47823 28070
rect 47857 28092 47860 28101
rect 47912 28092 47918 28144
rect 53208 28141 53236 28172
rect 53466 28160 53472 28212
rect 53524 28200 53530 28212
rect 53929 28203 53987 28209
rect 53929 28200 53941 28203
rect 53524 28172 53941 28200
rect 53524 28160 53530 28172
rect 53929 28169 53941 28172
rect 53975 28169 53987 28203
rect 53929 28163 53987 28169
rect 54665 28203 54723 28209
rect 54665 28169 54677 28203
rect 54711 28200 54723 28203
rect 55490 28200 55496 28212
rect 54711 28172 55496 28200
rect 54711 28169 54723 28172
rect 54665 28163 54723 28169
rect 55490 28160 55496 28172
rect 55548 28160 55554 28212
rect 51353 28135 51411 28141
rect 49344 28104 50200 28132
rect 47857 28067 47869 28092
rect 46716 28036 46761 28064
rect 47811 28061 47869 28067
rect 46716 28024 46722 28036
rect 48038 28024 48044 28076
rect 48096 28064 48102 28076
rect 48866 28064 48872 28076
rect 48096 28036 48872 28064
rect 48096 28024 48102 28036
rect 48866 28024 48872 28036
rect 48924 28024 48930 28076
rect 45741 27999 45799 28005
rect 45741 27965 45753 27999
rect 45787 27996 45799 27999
rect 45830 27996 45836 28008
rect 45787 27968 45836 27996
rect 45787 27965 45799 27968
rect 45741 27959 45799 27965
rect 45830 27956 45836 27968
rect 45888 27956 45894 28008
rect 47486 27956 47492 28008
rect 47544 27996 47550 28008
rect 49344 27996 49372 28104
rect 49421 28067 49479 28073
rect 49421 28033 49433 28067
rect 49467 28033 49479 28067
rect 49421 28027 49479 28033
rect 49605 28067 49663 28073
rect 49605 28033 49617 28067
rect 49651 28064 49663 28067
rect 49878 28064 49884 28076
rect 49651 28036 49884 28064
rect 49651 28033 49663 28036
rect 49605 28027 49663 28033
rect 47544 27968 49372 27996
rect 47544 27956 47550 27968
rect 43180 27900 44864 27928
rect 43916 27872 43944 27900
rect 45186 27888 45192 27940
rect 45244 27928 45250 27940
rect 48958 27928 48964 27940
rect 45244 27900 48964 27928
rect 45244 27888 45250 27900
rect 48958 27888 48964 27900
rect 49016 27928 49022 27940
rect 49436 27928 49464 28027
rect 49878 28024 49884 28036
rect 49936 28024 49942 28076
rect 50062 27996 50068 28008
rect 50023 27968 50068 27996
rect 50062 27956 50068 27968
rect 50120 27956 50126 28008
rect 49602 27928 49608 27940
rect 49016 27900 49608 27928
rect 49016 27888 49022 27900
rect 49602 27888 49608 27900
rect 49660 27888 49666 27940
rect 50172 27928 50200 28104
rect 51353 28101 51365 28135
rect 51399 28132 51411 28135
rect 53208 28135 53276 28141
rect 51399 28104 52960 28132
rect 53208 28104 53230 28135
rect 51399 28101 51411 28104
rect 51353 28095 51411 28101
rect 51074 28024 51080 28076
rect 51132 28064 51138 28076
rect 51537 28067 51595 28073
rect 51537 28064 51549 28067
rect 51132 28036 51549 28064
rect 51132 28024 51138 28036
rect 51537 28033 51549 28036
rect 51583 28033 51595 28067
rect 51537 28027 51595 28033
rect 51626 28024 51632 28076
rect 51684 28064 51690 28076
rect 51905 28067 51963 28073
rect 51684 28036 51729 28064
rect 51684 28024 51690 28036
rect 51905 28033 51917 28067
rect 51951 28033 51963 28067
rect 51905 28027 51963 28033
rect 52733 28067 52791 28073
rect 52733 28033 52745 28067
rect 52779 28064 52791 28067
rect 52822 28064 52828 28076
rect 52779 28036 52828 28064
rect 52779 28033 52791 28036
rect 52733 28027 52791 28033
rect 51350 27956 51356 28008
rect 51408 27996 51414 28008
rect 51920 27996 51948 28027
rect 52822 28024 52828 28036
rect 52880 28024 52886 28076
rect 52932 28064 52960 28104
rect 53218 28101 53230 28104
rect 53264 28101 53276 28135
rect 53218 28095 53276 28101
rect 53837 28067 53895 28073
rect 53837 28064 53849 28067
rect 52932 28036 53849 28064
rect 53837 28033 53849 28036
rect 53883 28033 53895 28067
rect 53837 28027 53895 28033
rect 54021 28067 54079 28073
rect 54021 28033 54033 28067
rect 54067 28033 54079 28067
rect 54478 28064 54484 28076
rect 54439 28036 54484 28064
rect 54021 28027 54079 28033
rect 51408 27968 51948 27996
rect 51408 27956 51414 27968
rect 52362 27956 52368 28008
rect 52420 27996 52426 28008
rect 53009 27999 53067 28005
rect 53009 27996 53021 27999
rect 52420 27968 53021 27996
rect 52420 27956 52426 27968
rect 53009 27965 53021 27968
rect 53055 27965 53067 27999
rect 53009 27959 53067 27965
rect 53098 27956 53104 28008
rect 53156 27996 53162 28008
rect 53156 27968 53201 27996
rect 53156 27956 53162 27968
rect 51813 27931 51871 27937
rect 51813 27928 51825 27931
rect 50172 27900 51825 27928
rect 51813 27897 51825 27900
rect 51859 27897 51871 27931
rect 51813 27891 51871 27897
rect 51902 27888 51908 27940
rect 51960 27928 51966 27940
rect 54036 27928 54064 28027
rect 54478 28024 54484 28036
rect 54536 28024 54542 28076
rect 54662 28064 54668 28076
rect 54623 28036 54668 28064
rect 54662 28024 54668 28036
rect 54720 28024 54726 28076
rect 56318 28024 56324 28076
rect 56376 28064 56382 28076
rect 58069 28067 58127 28073
rect 58069 28064 58081 28067
rect 56376 28036 58081 28064
rect 56376 28024 56382 28036
rect 58069 28033 58081 28036
rect 58115 28033 58127 28067
rect 58069 28027 58127 28033
rect 51960 27900 54064 27928
rect 51960 27888 51966 27900
rect 37884 27832 39436 27860
rect 41141 27863 41199 27869
rect 37884 27820 37890 27832
rect 41141 27829 41153 27863
rect 41187 27860 41199 27863
rect 43806 27860 43812 27872
rect 41187 27832 43812 27860
rect 41187 27829 41199 27832
rect 41141 27823 41199 27829
rect 43806 27820 43812 27832
rect 43864 27820 43870 27872
rect 43898 27820 43904 27872
rect 43956 27820 43962 27872
rect 45278 27820 45284 27872
rect 45336 27860 45342 27872
rect 46569 27863 46627 27869
rect 46569 27860 46581 27863
rect 45336 27832 46581 27860
rect 45336 27820 45342 27832
rect 46569 27829 46581 27832
rect 46615 27829 46627 27863
rect 47762 27860 47768 27872
rect 47723 27832 47768 27860
rect 46569 27823 46627 27829
rect 47762 27820 47768 27832
rect 47820 27820 47826 27872
rect 52454 27820 52460 27872
rect 52512 27860 52518 27872
rect 53098 27860 53104 27872
rect 52512 27832 53104 27860
rect 52512 27820 52518 27832
rect 53098 27820 53104 27832
rect 53156 27820 53162 27872
rect 53377 27863 53435 27869
rect 53377 27829 53389 27863
rect 53423 27860 53435 27863
rect 53650 27860 53656 27872
rect 53423 27832 53656 27860
rect 53423 27829 53435 27832
rect 53377 27823 53435 27829
rect 53650 27820 53656 27832
rect 53708 27820 53714 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 28810 27656 28816 27668
rect 28723 27628 28816 27656
rect 28810 27616 28816 27628
rect 28868 27656 28874 27668
rect 31662 27656 31668 27668
rect 28868 27628 31668 27656
rect 28868 27616 28874 27628
rect 31662 27616 31668 27628
rect 31720 27656 31726 27668
rect 31846 27656 31852 27668
rect 31720 27628 31852 27656
rect 31720 27616 31726 27628
rect 31846 27616 31852 27628
rect 31904 27616 31910 27668
rect 32677 27659 32735 27665
rect 32677 27656 32689 27659
rect 32140 27628 32689 27656
rect 28997 27591 29055 27597
rect 28997 27557 29009 27591
rect 29043 27588 29055 27591
rect 31570 27588 31576 27600
rect 29043 27560 31576 27588
rect 29043 27557 29055 27560
rect 28997 27551 29055 27557
rect 31570 27548 31576 27560
rect 31628 27548 31634 27600
rect 31754 27548 31760 27600
rect 31812 27588 31818 27600
rect 31812 27560 31892 27588
rect 31812 27548 31818 27560
rect 29270 27520 29276 27532
rect 28000 27492 29276 27520
rect 1946 27412 1952 27464
rect 2004 27452 2010 27464
rect 28000 27461 28028 27492
rect 29270 27480 29276 27492
rect 29328 27480 29334 27532
rect 30929 27523 30987 27529
rect 30929 27520 30941 27523
rect 29380 27492 30941 27520
rect 2225 27455 2283 27461
rect 2225 27452 2237 27455
rect 2004 27424 2237 27452
rect 2004 27412 2010 27424
rect 2225 27421 2237 27424
rect 2271 27421 2283 27455
rect 2225 27415 2283 27421
rect 27985 27455 28043 27461
rect 27985 27421 27997 27455
rect 28031 27421 28043 27455
rect 27985 27415 28043 27421
rect 28169 27455 28227 27461
rect 28169 27421 28181 27455
rect 28215 27452 28227 27455
rect 29086 27452 29092 27464
rect 28215 27424 29092 27452
rect 28215 27421 28227 27424
rect 28169 27415 28227 27421
rect 29086 27412 29092 27424
rect 29144 27412 29150 27464
rect 28629 27387 28687 27393
rect 28629 27353 28641 27387
rect 28675 27384 28687 27387
rect 28718 27384 28724 27396
rect 28675 27356 28724 27384
rect 28675 27353 28687 27356
rect 28629 27347 28687 27353
rect 28718 27344 28724 27356
rect 28776 27344 28782 27396
rect 28845 27387 28903 27393
rect 28845 27384 28857 27387
rect 28828 27353 28857 27384
rect 28891 27384 28903 27387
rect 28891 27356 29132 27384
rect 28891 27353 28903 27356
rect 28828 27347 28903 27353
rect 28169 27319 28227 27325
rect 28169 27285 28181 27319
rect 28215 27316 28227 27319
rect 28828 27316 28856 27347
rect 28215 27288 28856 27316
rect 29104 27316 29132 27356
rect 29380 27316 29408 27492
rect 30929 27489 30941 27492
rect 30975 27489 30987 27523
rect 30929 27483 30987 27489
rect 31294 27480 31300 27532
rect 31352 27520 31358 27532
rect 31864 27529 31892 27560
rect 31657 27523 31715 27529
rect 31657 27520 31669 27523
rect 31352 27492 31669 27520
rect 31352 27480 31358 27492
rect 31657 27489 31669 27492
rect 31703 27489 31715 27523
rect 31657 27483 31715 27489
rect 31849 27523 31907 27529
rect 31849 27489 31861 27523
rect 31895 27489 31907 27523
rect 31849 27483 31907 27489
rect 31942 27523 32000 27529
rect 31942 27489 31954 27523
rect 31988 27520 32000 27523
rect 32030 27520 32036 27532
rect 31988 27492 32036 27520
rect 31988 27489 32000 27492
rect 31942 27483 32000 27489
rect 32030 27480 32036 27492
rect 32088 27480 32094 27532
rect 30466 27452 30472 27464
rect 30427 27424 30472 27452
rect 30466 27412 30472 27424
rect 30524 27412 30530 27464
rect 30561 27455 30619 27461
rect 30561 27421 30573 27455
rect 30607 27452 30619 27455
rect 30742 27452 30748 27464
rect 30607 27424 30748 27452
rect 30607 27421 30619 27424
rect 30561 27415 30619 27421
rect 30742 27412 30748 27424
rect 30800 27412 30806 27464
rect 30837 27455 30895 27461
rect 30837 27421 30849 27455
rect 30883 27452 30895 27455
rect 31478 27452 31484 27464
rect 30883 27424 31484 27452
rect 30883 27421 30895 27424
rect 30837 27415 30895 27421
rect 29822 27384 29828 27396
rect 29783 27356 29828 27384
rect 29822 27344 29828 27356
rect 29880 27344 29886 27396
rect 30282 27344 30288 27396
rect 30340 27384 30346 27396
rect 30852 27384 30880 27415
rect 31478 27412 31484 27424
rect 31536 27412 31542 27464
rect 31570 27412 31576 27464
rect 31628 27452 31634 27464
rect 31757 27455 31815 27461
rect 31757 27452 31769 27455
rect 31628 27424 31769 27452
rect 31628 27412 31634 27424
rect 31757 27421 31769 27424
rect 31803 27454 31815 27455
rect 31803 27452 31984 27454
rect 32140 27452 32168 27628
rect 32677 27625 32689 27628
rect 32723 27656 32735 27659
rect 33042 27656 33048 27668
rect 32723 27628 33048 27656
rect 32723 27625 32735 27628
rect 32677 27619 32735 27625
rect 33042 27616 33048 27628
rect 33100 27616 33106 27668
rect 36354 27616 36360 27668
rect 36412 27656 36418 27668
rect 37093 27659 37151 27665
rect 37093 27656 37105 27659
rect 36412 27628 37105 27656
rect 36412 27616 36418 27628
rect 37093 27625 37105 27628
rect 37139 27625 37151 27659
rect 37093 27619 37151 27625
rect 37182 27616 37188 27668
rect 37240 27656 37246 27668
rect 37921 27659 37979 27665
rect 37921 27656 37933 27659
rect 37240 27628 37933 27656
rect 37240 27616 37246 27628
rect 37921 27625 37933 27628
rect 37967 27625 37979 27659
rect 37921 27619 37979 27625
rect 38010 27616 38016 27668
rect 38068 27656 38074 27668
rect 38105 27659 38163 27665
rect 38105 27656 38117 27659
rect 38068 27628 38117 27656
rect 38068 27616 38074 27628
rect 38105 27625 38117 27628
rect 38151 27625 38163 27659
rect 38105 27619 38163 27625
rect 38194 27616 38200 27668
rect 38252 27656 38258 27668
rect 38749 27659 38807 27665
rect 38749 27656 38761 27659
rect 38252 27628 38761 27656
rect 38252 27616 38258 27628
rect 38749 27625 38761 27628
rect 38795 27625 38807 27659
rect 38749 27619 38807 27625
rect 41046 27616 41052 27668
rect 41104 27656 41110 27668
rect 41690 27656 41696 27668
rect 41104 27628 41696 27656
rect 41104 27616 41110 27628
rect 41690 27616 41696 27628
rect 41748 27616 41754 27668
rect 43714 27616 43720 27668
rect 43772 27656 43778 27668
rect 43993 27659 44051 27665
rect 43993 27656 44005 27659
rect 43772 27628 44005 27656
rect 43772 27616 43778 27628
rect 43993 27625 44005 27628
rect 44039 27625 44051 27659
rect 43993 27619 44051 27625
rect 44652 27628 45140 27656
rect 32858 27548 32864 27600
rect 32916 27588 32922 27600
rect 33413 27591 33471 27597
rect 33413 27588 33425 27591
rect 32916 27560 33425 27588
rect 32916 27548 32922 27560
rect 33413 27557 33425 27560
rect 33459 27557 33471 27591
rect 36170 27588 36176 27600
rect 36083 27560 36176 27588
rect 33413 27551 33471 27557
rect 36170 27548 36176 27560
rect 36228 27588 36234 27600
rect 40681 27591 40739 27597
rect 36228 27560 38654 27588
rect 36228 27548 36234 27560
rect 36188 27461 36216 27548
rect 36265 27523 36323 27529
rect 36265 27489 36277 27523
rect 36311 27520 36323 27523
rect 36817 27523 36875 27529
rect 36817 27520 36829 27523
rect 36311 27492 36829 27520
rect 36311 27489 36323 27492
rect 36265 27483 36323 27489
rect 36817 27489 36829 27492
rect 36863 27520 36875 27523
rect 38010 27520 38016 27532
rect 36863 27492 38016 27520
rect 36863 27489 36875 27492
rect 36817 27483 36875 27489
rect 38010 27480 38016 27492
rect 38068 27480 38074 27532
rect 38626 27520 38654 27560
rect 40681 27557 40693 27591
rect 40727 27588 40739 27591
rect 44652 27588 44680 27628
rect 40727 27560 44680 27588
rect 40727 27557 40739 27560
rect 40681 27551 40739 27557
rect 44726 27548 44732 27600
rect 44784 27588 44790 27600
rect 45005 27591 45063 27597
rect 45005 27588 45017 27591
rect 44784 27560 45017 27588
rect 44784 27548 44790 27560
rect 45005 27557 45017 27560
rect 45051 27557 45063 27591
rect 45112 27588 45140 27628
rect 45186 27616 45192 27668
rect 45244 27656 45250 27668
rect 45922 27656 45928 27668
rect 45244 27628 45928 27656
rect 45244 27616 45250 27628
rect 45922 27616 45928 27628
rect 45980 27656 45986 27668
rect 46017 27659 46075 27665
rect 46017 27656 46029 27659
rect 45980 27628 46029 27656
rect 45980 27616 45986 27628
rect 46017 27625 46029 27628
rect 46063 27625 46075 27659
rect 46382 27656 46388 27668
rect 46343 27628 46388 27656
rect 46017 27619 46075 27625
rect 46382 27616 46388 27628
rect 46440 27616 46446 27668
rect 47397 27659 47455 27665
rect 47397 27625 47409 27659
rect 47443 27656 47455 27659
rect 47762 27656 47768 27668
rect 47443 27628 47768 27656
rect 47443 27625 47455 27628
rect 47397 27619 47455 27625
rect 47762 27616 47768 27628
rect 47820 27616 47826 27668
rect 47854 27616 47860 27668
rect 47912 27656 47918 27668
rect 47949 27659 48007 27665
rect 47949 27656 47961 27659
rect 47912 27628 47961 27656
rect 47912 27616 47918 27628
rect 47949 27625 47961 27628
rect 47995 27625 48007 27659
rect 52914 27656 52920 27668
rect 52875 27628 52920 27656
rect 47949 27619 48007 27625
rect 52914 27616 52920 27628
rect 52972 27616 52978 27668
rect 48866 27588 48872 27600
rect 45112 27560 48872 27588
rect 45005 27551 45063 27557
rect 48866 27548 48872 27560
rect 48924 27588 48930 27600
rect 49605 27591 49663 27597
rect 48924 27560 49372 27588
rect 48924 27548 48930 27560
rect 47489 27523 47547 27529
rect 38626 27492 46060 27520
rect 33321 27455 33379 27461
rect 33321 27452 33333 27455
rect 31803 27426 32168 27452
rect 31803 27421 31815 27426
rect 31956 27424 32168 27426
rect 32324 27424 33333 27452
rect 31757 27415 31815 27421
rect 30340 27356 30880 27384
rect 31496 27384 31524 27412
rect 31938 27384 31944 27396
rect 31496 27356 31944 27384
rect 30340 27344 30346 27356
rect 31938 27344 31944 27356
rect 31996 27384 32002 27396
rect 32324 27384 32352 27424
rect 33321 27421 33333 27424
rect 33367 27421 33379 27455
rect 33321 27415 33379 27421
rect 33505 27455 33563 27461
rect 33505 27421 33517 27455
rect 33551 27421 33563 27455
rect 33505 27415 33563 27421
rect 36173 27455 36231 27461
rect 36173 27421 36185 27455
rect 36219 27421 36231 27455
rect 36354 27452 36360 27464
rect 36315 27424 36360 27452
rect 36173 27415 36231 27421
rect 32490 27384 32496 27396
rect 31996 27356 32352 27384
rect 32451 27356 32496 27384
rect 31996 27344 32002 27356
rect 32490 27344 32496 27356
rect 32548 27384 32554 27396
rect 33520 27384 33548 27415
rect 36354 27412 36360 27424
rect 36412 27412 36418 27464
rect 37090 27452 37096 27464
rect 37051 27424 37096 27452
rect 37090 27412 37096 27424
rect 37148 27412 37154 27464
rect 37277 27455 37335 27461
rect 37277 27421 37289 27455
rect 37323 27452 37335 27455
rect 37366 27452 37372 27464
rect 37323 27424 37372 27452
rect 37323 27421 37335 27424
rect 37277 27415 37335 27421
rect 37366 27412 37372 27424
rect 37424 27452 37430 27464
rect 37642 27452 37648 27464
rect 37424 27424 37648 27452
rect 37424 27412 37430 27424
rect 37642 27412 37648 27424
rect 37700 27412 37706 27464
rect 37826 27412 37832 27464
rect 37884 27452 37890 27464
rect 38565 27455 38623 27461
rect 38565 27452 38577 27455
rect 37884 27424 38577 27452
rect 37884 27412 37890 27424
rect 38565 27421 38577 27424
rect 38611 27421 38623 27455
rect 38565 27415 38623 27421
rect 41506 27412 41512 27464
rect 41564 27452 41570 27464
rect 41782 27452 41788 27464
rect 41564 27424 41609 27452
rect 41743 27424 41788 27452
rect 41564 27412 41570 27424
rect 41782 27412 41788 27424
rect 41840 27412 41846 27464
rect 42334 27452 42340 27464
rect 42295 27424 42340 27452
rect 42334 27412 42340 27424
rect 42392 27412 42398 27464
rect 43625 27455 43683 27461
rect 43625 27421 43637 27455
rect 43671 27452 43683 27455
rect 43898 27452 43904 27464
rect 43671 27424 43904 27452
rect 43671 27421 43683 27424
rect 43625 27415 43683 27421
rect 43898 27412 43904 27424
rect 43956 27412 43962 27464
rect 45186 27452 45192 27464
rect 45147 27424 45192 27452
rect 45186 27412 45192 27424
rect 45244 27412 45250 27464
rect 45465 27455 45523 27461
rect 45465 27421 45477 27455
rect 45511 27452 45523 27455
rect 45738 27452 45744 27464
rect 45511 27424 45744 27452
rect 45511 27421 45523 27424
rect 45465 27415 45523 27421
rect 45738 27412 45744 27424
rect 45796 27412 45802 27464
rect 45922 27452 45928 27464
rect 45883 27424 45928 27452
rect 45922 27412 45928 27424
rect 45980 27412 45986 27464
rect 32548 27356 33548 27384
rect 37737 27387 37795 27393
rect 32548 27344 32554 27356
rect 37737 27353 37749 27387
rect 37783 27353 37795 27387
rect 37737 27347 37795 27353
rect 37953 27387 38011 27393
rect 37953 27353 37965 27387
rect 37999 27384 38011 27387
rect 38286 27384 38292 27396
rect 37999 27356 38292 27384
rect 37999 27353 38011 27356
rect 37953 27347 38011 27353
rect 29104 27288 29408 27316
rect 28215 27285 28227 27288
rect 28169 27279 28227 27285
rect 30374 27276 30380 27328
rect 30432 27316 30438 27328
rect 31481 27319 31539 27325
rect 31481 27316 31493 27319
rect 30432 27288 31493 27316
rect 30432 27276 30438 27288
rect 31481 27285 31493 27288
rect 31527 27285 31539 27319
rect 31481 27279 31539 27285
rect 32122 27276 32128 27328
rect 32180 27316 32186 27328
rect 32693 27319 32751 27325
rect 32693 27316 32705 27319
rect 32180 27288 32705 27316
rect 32180 27276 32186 27288
rect 32693 27285 32705 27288
rect 32739 27285 32751 27319
rect 32858 27316 32864 27328
rect 32819 27288 32864 27316
rect 32693 27279 32751 27285
rect 32858 27276 32864 27288
rect 32916 27276 32922 27328
rect 36722 27276 36728 27328
rect 36780 27316 36786 27328
rect 37752 27316 37780 27347
rect 38286 27344 38292 27356
rect 38344 27344 38350 27396
rect 40497 27387 40555 27393
rect 40497 27384 40509 27387
rect 38396 27356 40509 27384
rect 38396 27316 38424 27356
rect 40497 27353 40509 27356
rect 40543 27353 40555 27387
rect 40497 27347 40555 27353
rect 41690 27344 41696 27396
rect 41748 27384 41754 27396
rect 42521 27387 42579 27393
rect 41748 27356 41793 27384
rect 41748 27344 41754 27356
rect 42521 27353 42533 27387
rect 42567 27384 42579 27387
rect 42794 27384 42800 27396
rect 42567 27356 42800 27384
rect 42567 27353 42579 27356
rect 42521 27347 42579 27353
rect 42794 27344 42800 27356
rect 42852 27384 42858 27396
rect 43254 27384 43260 27396
rect 42852 27356 43260 27384
rect 42852 27344 42858 27356
rect 43254 27344 43260 27356
rect 43312 27384 43318 27396
rect 43809 27387 43867 27393
rect 43809 27384 43821 27387
rect 43312 27356 43821 27384
rect 43312 27344 43318 27356
rect 43809 27353 43821 27356
rect 43855 27353 43867 27387
rect 43809 27347 43867 27353
rect 36780 27288 38424 27316
rect 36780 27276 36786 27288
rect 39482 27276 39488 27328
rect 39540 27316 39546 27328
rect 40586 27316 40592 27328
rect 39540 27288 40592 27316
rect 39540 27276 39546 27288
rect 40586 27276 40592 27288
rect 40644 27276 40650 27328
rect 41325 27319 41383 27325
rect 41325 27285 41337 27319
rect 41371 27316 41383 27319
rect 42334 27316 42340 27328
rect 41371 27288 42340 27316
rect 41371 27285 41383 27288
rect 41325 27279 41383 27285
rect 42334 27276 42340 27288
rect 42392 27276 42398 27328
rect 45370 27276 45376 27328
rect 45428 27316 45434 27328
rect 45922 27316 45928 27328
rect 45428 27288 45928 27316
rect 45428 27276 45434 27288
rect 45922 27276 45928 27288
rect 45980 27276 45986 27328
rect 46032 27316 46060 27492
rect 47489 27489 47501 27523
rect 47535 27520 47547 27523
rect 47670 27520 47676 27532
rect 47535 27492 47676 27520
rect 47535 27489 47547 27492
rect 47489 27483 47547 27489
rect 47670 27480 47676 27492
rect 47728 27480 47734 27532
rect 49344 27520 49372 27560
rect 49605 27557 49617 27591
rect 49651 27588 49663 27591
rect 56962 27588 56968 27600
rect 49651 27560 51074 27588
rect 56923 27560 56968 27588
rect 49651 27557 49663 27560
rect 49605 27551 49663 27557
rect 47872 27492 48544 27520
rect 46290 27412 46296 27464
rect 46348 27452 46354 27464
rect 47213 27455 47271 27461
rect 47213 27452 47225 27455
rect 46348 27424 47225 27452
rect 46348 27412 46354 27424
rect 47213 27421 47225 27424
rect 47259 27421 47271 27455
rect 47213 27415 47271 27421
rect 47228 27384 47256 27415
rect 47302 27412 47308 27464
rect 47360 27452 47366 27464
rect 47872 27452 47900 27492
rect 48130 27452 48136 27464
rect 47360 27424 47900 27452
rect 48091 27424 48136 27452
rect 47360 27412 47366 27424
rect 48130 27412 48136 27424
rect 48188 27412 48194 27464
rect 48225 27455 48283 27461
rect 48225 27421 48237 27455
rect 48271 27452 48283 27455
rect 48314 27452 48320 27464
rect 48271 27424 48320 27452
rect 48271 27421 48283 27424
rect 48225 27415 48283 27421
rect 48314 27412 48320 27424
rect 48372 27412 48378 27464
rect 48516 27461 48544 27492
rect 49344 27492 49648 27520
rect 49344 27461 49372 27492
rect 48409 27455 48467 27461
rect 48409 27421 48421 27455
rect 48455 27421 48467 27455
rect 48409 27415 48467 27421
rect 48501 27455 48559 27461
rect 48501 27421 48513 27455
rect 48547 27421 48559 27455
rect 48501 27415 48559 27421
rect 49053 27455 49111 27461
rect 49053 27421 49065 27455
rect 49099 27421 49111 27455
rect 49053 27415 49111 27421
rect 49329 27455 49387 27461
rect 49329 27421 49341 27455
rect 49375 27421 49387 27455
rect 49329 27415 49387 27421
rect 48424 27384 48452 27415
rect 47228 27356 48452 27384
rect 49068 27316 49096 27415
rect 49418 27412 49424 27464
rect 49476 27452 49482 27464
rect 49620 27452 49648 27492
rect 49878 27480 49884 27532
rect 49936 27520 49942 27532
rect 50433 27523 50491 27529
rect 50433 27520 50445 27523
rect 49936 27492 50445 27520
rect 49936 27480 49942 27492
rect 50433 27489 50445 27492
rect 50479 27489 50491 27523
rect 51046 27520 51074 27560
rect 56962 27548 56968 27560
rect 57020 27548 57026 27600
rect 53006 27520 53012 27532
rect 51046 27492 53012 27520
rect 50433 27483 50491 27489
rect 50157 27455 50215 27461
rect 50157 27452 50169 27455
rect 49476 27424 49521 27452
rect 49620 27424 50169 27452
rect 49476 27412 49482 27424
rect 50157 27421 50169 27424
rect 50203 27421 50215 27455
rect 51442 27452 51448 27464
rect 51403 27424 51448 27452
rect 50157 27415 50215 27421
rect 51442 27412 51448 27424
rect 51500 27412 51506 27464
rect 51721 27455 51779 27461
rect 51721 27421 51733 27455
rect 51767 27452 51779 27455
rect 52362 27452 52368 27464
rect 51767 27424 52368 27452
rect 51767 27421 51779 27424
rect 51721 27415 51779 27421
rect 49234 27384 49240 27396
rect 49195 27356 49240 27384
rect 49234 27344 49240 27356
rect 49292 27344 49298 27396
rect 49602 27344 49608 27396
rect 49660 27384 49666 27396
rect 50798 27384 50804 27396
rect 49660 27356 50804 27384
rect 49660 27344 49666 27356
rect 50798 27344 50804 27356
rect 50856 27384 50862 27396
rect 50856 27356 51074 27384
rect 50856 27344 50862 27356
rect 50154 27316 50160 27328
rect 46032 27288 50160 27316
rect 50154 27276 50160 27288
rect 50212 27276 50218 27328
rect 51046 27316 51074 27356
rect 51166 27344 51172 27396
rect 51224 27384 51230 27396
rect 51736 27384 51764 27415
rect 52362 27412 52368 27424
rect 52420 27412 52426 27464
rect 52748 27461 52776 27492
rect 53006 27480 53012 27492
rect 53064 27480 53070 27532
rect 53561 27523 53619 27529
rect 53561 27489 53573 27523
rect 53607 27520 53619 27523
rect 54478 27520 54484 27532
rect 53607 27492 54484 27520
rect 53607 27489 53619 27492
rect 53561 27483 53619 27489
rect 54478 27480 54484 27492
rect 54536 27480 54542 27532
rect 52733 27455 52791 27461
rect 52733 27421 52745 27455
rect 52779 27421 52791 27455
rect 52733 27415 52791 27421
rect 53190 27412 53196 27464
rect 53248 27452 53254 27464
rect 53469 27455 53527 27461
rect 53469 27452 53481 27455
rect 53248 27424 53481 27452
rect 53248 27412 53254 27424
rect 53469 27421 53481 27424
rect 53515 27421 53527 27455
rect 53650 27452 53656 27464
rect 53611 27424 53656 27452
rect 53469 27415 53527 27421
rect 53650 27412 53656 27424
rect 53708 27412 53714 27464
rect 56778 27412 56784 27464
rect 56836 27452 56842 27464
rect 56873 27455 56931 27461
rect 56873 27452 56885 27455
rect 56836 27424 56885 27452
rect 56836 27412 56842 27424
rect 56873 27421 56885 27424
rect 56919 27421 56931 27455
rect 56873 27415 56931 27421
rect 51224 27356 51764 27384
rect 51224 27344 51230 27356
rect 51534 27316 51540 27328
rect 51046 27288 51540 27316
rect 51534 27276 51540 27288
rect 51592 27276 51598 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 8478 27072 8484 27124
rect 8536 27112 8542 27124
rect 29822 27112 29828 27124
rect 8536 27084 29828 27112
rect 8536 27072 8542 27084
rect 29822 27072 29828 27084
rect 29880 27072 29886 27124
rect 30742 27072 30748 27124
rect 30800 27112 30806 27124
rect 31478 27112 31484 27124
rect 30800 27084 31484 27112
rect 30800 27072 30806 27084
rect 31478 27072 31484 27084
rect 31536 27112 31542 27124
rect 32585 27115 32643 27121
rect 32585 27112 32597 27115
rect 31536 27084 32597 27112
rect 31536 27072 31542 27084
rect 32585 27081 32597 27084
rect 32631 27081 32643 27115
rect 37734 27112 37740 27124
rect 37695 27084 37740 27112
rect 32585 27075 32643 27081
rect 37734 27072 37740 27084
rect 37792 27072 37798 27124
rect 41506 27112 41512 27124
rect 41156 27084 41512 27112
rect 28721 27047 28779 27053
rect 28721 27013 28733 27047
rect 28767 27044 28779 27047
rect 30466 27044 30472 27056
rect 28767 27016 30472 27044
rect 28767 27013 28779 27016
rect 28721 27007 28779 27013
rect 30466 27004 30472 27016
rect 30524 27004 30530 27056
rect 31294 27044 31300 27056
rect 31036 27016 31300 27044
rect 1946 26976 1952 26988
rect 1907 26948 1952 26976
rect 1946 26936 1952 26948
rect 2004 26936 2010 26988
rect 8754 26976 8760 26988
rect 8715 26948 8760 26976
rect 8754 26936 8760 26948
rect 8812 26936 8818 26988
rect 28629 26979 28687 26985
rect 28629 26945 28641 26979
rect 28675 26945 28687 26979
rect 28629 26939 28687 26945
rect 28813 26979 28871 26985
rect 28813 26945 28825 26979
rect 28859 26945 28871 26979
rect 28813 26939 28871 26945
rect 29273 26979 29331 26985
rect 29273 26945 29285 26979
rect 29319 26945 29331 26979
rect 29273 26939 29331 26945
rect 29457 26979 29515 26985
rect 29457 26945 29469 26979
rect 29503 26976 29515 26979
rect 29546 26976 29552 26988
rect 29503 26948 29552 26976
rect 29503 26945 29515 26948
rect 29457 26939 29515 26945
rect 2133 26911 2191 26917
rect 2133 26877 2145 26911
rect 2179 26908 2191 26911
rect 2498 26908 2504 26920
rect 2179 26880 2504 26908
rect 2179 26877 2191 26880
rect 2133 26871 2191 26877
rect 2498 26868 2504 26880
rect 2556 26868 2562 26920
rect 2774 26908 2780 26920
rect 2735 26880 2780 26908
rect 2774 26868 2780 26880
rect 2832 26868 2838 26920
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 9033 26911 9091 26917
rect 9033 26908 9045 26911
rect 8628 26880 9045 26908
rect 8628 26868 8634 26880
rect 9033 26877 9045 26880
rect 9079 26877 9091 26911
rect 9033 26871 9091 26877
rect 28644 26772 28672 26939
rect 28828 26852 28856 26939
rect 28994 26908 29000 26920
rect 28966 26868 29000 26908
rect 29052 26868 29058 26920
rect 28810 26800 28816 26852
rect 28868 26800 28874 26852
rect 28966 26772 28994 26868
rect 29288 26840 29316 26939
rect 29546 26936 29552 26948
rect 29604 26936 29610 26988
rect 29730 26936 29736 26988
rect 29788 26976 29794 26988
rect 31036 26976 31064 27016
rect 31294 27004 31300 27016
rect 31352 27044 31358 27056
rect 32122 27044 32128 27056
rect 31352 27016 31432 27044
rect 32083 27016 32128 27044
rect 31352 27004 31358 27016
rect 29788 26948 31064 26976
rect 29788 26936 29794 26948
rect 31110 26936 31116 26988
rect 31168 26976 31174 26988
rect 31404 26985 31432 27016
rect 32122 27004 32128 27016
rect 32180 27004 32186 27056
rect 36814 27044 36820 27056
rect 36556 27016 36820 27044
rect 36556 26985 36584 27016
rect 36814 27004 36820 27016
rect 36872 27044 36878 27056
rect 36872 27016 37596 27044
rect 36872 27004 36878 27016
rect 31389 26979 31447 26985
rect 31168 26948 31340 26976
rect 31168 26936 31174 26948
rect 31312 26920 31340 26948
rect 31389 26945 31401 26979
rect 31435 26945 31447 26979
rect 31389 26939 31447 26945
rect 36541 26979 36599 26985
rect 36541 26945 36553 26979
rect 36587 26945 36599 26979
rect 36722 26976 36728 26988
rect 36683 26948 36728 26976
rect 36541 26939 36599 26945
rect 36722 26936 36728 26948
rect 36780 26936 36786 26988
rect 37568 26985 37596 27016
rect 38838 27004 38844 27056
rect 38896 27044 38902 27056
rect 39485 27047 39543 27053
rect 39485 27044 39497 27047
rect 38896 27016 39497 27044
rect 38896 27004 38902 27016
rect 39485 27013 39497 27016
rect 39531 27013 39543 27047
rect 40494 27044 40500 27056
rect 39485 27007 39543 27013
rect 40144 27016 40500 27044
rect 37553 26979 37611 26985
rect 37553 26945 37565 26979
rect 37599 26945 37611 26979
rect 37826 26976 37832 26988
rect 37739 26948 37832 26976
rect 37553 26939 37611 26945
rect 37826 26936 37832 26948
rect 37884 26976 37890 26988
rect 38378 26976 38384 26988
rect 37884 26948 38384 26976
rect 37884 26936 37890 26948
rect 38378 26936 38384 26948
rect 38436 26936 38442 26988
rect 40144 26985 40172 27016
rect 40494 27004 40500 27016
rect 40552 27004 40558 27056
rect 40129 26979 40187 26985
rect 40129 26976 40141 26979
rect 38948 26948 40141 26976
rect 29638 26868 29644 26920
rect 29696 26908 29702 26920
rect 29917 26911 29975 26917
rect 29917 26908 29929 26911
rect 29696 26880 29929 26908
rect 29696 26868 29702 26880
rect 29917 26877 29929 26880
rect 29963 26908 29975 26911
rect 30006 26908 30012 26920
rect 29963 26880 30012 26908
rect 29963 26877 29975 26880
rect 29917 26871 29975 26877
rect 30006 26868 30012 26880
rect 30064 26868 30070 26920
rect 30193 26911 30251 26917
rect 30193 26877 30205 26911
rect 30239 26908 30251 26911
rect 30926 26908 30932 26920
rect 30239 26880 30932 26908
rect 30239 26877 30251 26880
rect 30193 26871 30251 26877
rect 30926 26868 30932 26880
rect 30984 26908 30990 26920
rect 31202 26908 31208 26920
rect 30984 26880 31208 26908
rect 30984 26868 30990 26880
rect 31202 26868 31208 26880
rect 31260 26868 31266 26920
rect 31294 26868 31300 26920
rect 31352 26908 31358 26920
rect 32490 26908 32496 26920
rect 31352 26880 32496 26908
rect 31352 26868 31358 26880
rect 32490 26868 32496 26880
rect 32548 26868 32554 26920
rect 36633 26911 36691 26917
rect 36633 26877 36645 26911
rect 36679 26908 36691 26911
rect 37642 26908 37648 26920
rect 36679 26880 37648 26908
rect 36679 26877 36691 26880
rect 36633 26871 36691 26877
rect 37642 26868 37648 26880
rect 37700 26868 37706 26920
rect 30834 26840 30840 26852
rect 29288 26812 30840 26840
rect 30834 26800 30840 26812
rect 30892 26840 30898 26852
rect 31573 26843 31631 26849
rect 31573 26840 31585 26843
rect 30892 26812 31585 26840
rect 30892 26800 30898 26812
rect 31573 26809 31585 26812
rect 31619 26809 31631 26843
rect 31573 26803 31631 26809
rect 32214 26800 32220 26852
rect 32272 26840 32278 26852
rect 32401 26843 32459 26849
rect 32401 26840 32413 26843
rect 32272 26812 32413 26840
rect 32272 26800 32278 26812
rect 32401 26809 32413 26812
rect 32447 26809 32459 26843
rect 32401 26803 32459 26809
rect 36538 26800 36544 26852
rect 36596 26840 36602 26852
rect 38948 26840 38976 26948
rect 40129 26945 40141 26948
rect 40175 26945 40187 26979
rect 40129 26939 40187 26945
rect 40313 26979 40371 26985
rect 40313 26945 40325 26979
rect 40359 26976 40371 26979
rect 40678 26976 40684 26988
rect 40359 26948 40684 26976
rect 40359 26945 40371 26948
rect 40313 26939 40371 26945
rect 40678 26936 40684 26948
rect 40736 26936 40742 26988
rect 40865 26979 40923 26985
rect 40865 26945 40877 26979
rect 40911 26976 40923 26979
rect 41046 26976 41052 26988
rect 40911 26948 41052 26976
rect 40911 26945 40923 26948
rect 40865 26939 40923 26945
rect 41046 26936 41052 26948
rect 41104 26936 41110 26988
rect 41156 26985 41184 27084
rect 41506 27072 41512 27084
rect 41564 27072 41570 27124
rect 44634 27072 44640 27124
rect 44692 27112 44698 27124
rect 46385 27115 46443 27121
rect 46385 27112 46397 27115
rect 44692 27084 46397 27112
rect 44692 27072 44698 27084
rect 46385 27081 46397 27084
rect 46431 27081 46443 27115
rect 46385 27075 46443 27081
rect 48130 27072 48136 27124
rect 48188 27112 48194 27124
rect 49237 27115 49295 27121
rect 49237 27112 49249 27115
rect 48188 27084 49249 27112
rect 48188 27072 48194 27084
rect 49237 27081 49249 27084
rect 49283 27081 49295 27115
rect 49237 27075 49295 27081
rect 49326 27072 49332 27124
rect 49384 27112 49390 27124
rect 51350 27112 51356 27124
rect 49384 27084 51356 27112
rect 49384 27072 49390 27084
rect 51350 27072 51356 27084
rect 51408 27072 51414 27124
rect 51534 27112 51540 27124
rect 51495 27084 51540 27112
rect 51534 27072 51540 27084
rect 51592 27072 51598 27124
rect 51813 27115 51871 27121
rect 51813 27081 51825 27115
rect 51859 27112 51871 27115
rect 51902 27112 51908 27124
rect 51859 27084 51908 27112
rect 51859 27081 51871 27084
rect 51813 27075 51871 27081
rect 51902 27072 51908 27084
rect 51960 27072 51966 27124
rect 55950 27072 55956 27124
rect 56008 27112 56014 27124
rect 57057 27115 57115 27121
rect 57057 27112 57069 27115
rect 56008 27084 57069 27112
rect 56008 27072 56014 27084
rect 57057 27081 57069 27084
rect 57103 27081 57115 27115
rect 57057 27075 57115 27081
rect 41230 27004 41236 27056
rect 41288 27044 41294 27056
rect 41288 27016 41333 27044
rect 41288 27004 41294 27016
rect 42334 27004 42340 27056
rect 42392 27044 42398 27056
rect 47302 27044 47308 27056
rect 42392 27016 47308 27044
rect 42392 27004 42398 27016
rect 41141 26979 41199 26985
rect 41141 26945 41153 26979
rect 41187 26945 41199 26979
rect 41141 26939 41199 26945
rect 41417 26979 41475 26985
rect 41417 26945 41429 26979
rect 41463 26976 41475 26979
rect 42794 26976 42800 26988
rect 41463 26948 42800 26976
rect 41463 26945 41475 26948
rect 41417 26939 41475 26945
rect 42794 26936 42800 26948
rect 42852 26936 42858 26988
rect 43714 26976 43720 26988
rect 43675 26948 43720 26976
rect 43714 26936 43720 26948
rect 43772 26936 43778 26988
rect 43901 26979 43959 26985
rect 43901 26945 43913 26979
rect 43947 26945 43959 26979
rect 46290 26976 46296 26988
rect 46251 26948 46296 26976
rect 43901 26939 43959 26945
rect 40218 26868 40224 26920
rect 40276 26908 40282 26920
rect 41693 26911 41751 26917
rect 41693 26908 41705 26911
rect 40276 26880 41705 26908
rect 40276 26868 40282 26880
rect 41693 26877 41705 26880
rect 41739 26877 41751 26911
rect 41693 26871 41751 26877
rect 43530 26868 43536 26920
rect 43588 26908 43594 26920
rect 43916 26908 43944 26939
rect 46290 26936 46296 26948
rect 46348 26936 46354 26988
rect 46768 26985 46796 27016
rect 47302 27004 47308 27016
rect 47360 27004 47366 27056
rect 48869 27047 48927 27053
rect 48869 27013 48881 27047
rect 48915 27044 48927 27047
rect 48958 27044 48964 27056
rect 48915 27016 48964 27044
rect 48915 27013 48927 27016
rect 48869 27007 48927 27013
rect 48958 27004 48964 27016
rect 49016 27004 49022 27056
rect 49053 27047 49111 27053
rect 49053 27013 49065 27047
rect 49099 27044 49111 27047
rect 49878 27044 49884 27056
rect 49099 27016 49884 27044
rect 49099 27013 49111 27016
rect 49053 27007 49111 27013
rect 49878 27004 49884 27016
rect 49936 27004 49942 27056
rect 51077 27047 51135 27053
rect 51077 27013 51089 27047
rect 51123 27044 51135 27047
rect 51626 27044 51632 27056
rect 51123 27016 51632 27044
rect 51123 27013 51135 27016
rect 51077 27007 51135 27013
rect 51626 27004 51632 27016
rect 51684 27004 51690 27056
rect 46753 26979 46811 26985
rect 46753 26945 46765 26979
rect 46799 26945 46811 26979
rect 48038 26976 48044 26988
rect 47999 26948 48044 26976
rect 46753 26939 46811 26945
rect 48038 26936 48044 26948
rect 48096 26936 48102 26988
rect 56594 26976 56600 26988
rect 49160 26948 56600 26976
rect 43588 26880 43944 26908
rect 43588 26868 43594 26880
rect 47118 26868 47124 26920
rect 47176 26908 47182 26920
rect 49160 26908 49188 26948
rect 56594 26936 56600 26948
rect 56652 26976 56658 26988
rect 56873 26979 56931 26985
rect 56873 26976 56885 26979
rect 56652 26948 56885 26976
rect 56652 26936 56658 26948
rect 56873 26945 56885 26948
rect 56919 26945 56931 26979
rect 56873 26939 56931 26945
rect 49694 26908 49700 26920
rect 47176 26880 49188 26908
rect 49655 26880 49700 26908
rect 47176 26868 47182 26880
rect 49694 26868 49700 26880
rect 49752 26868 49758 26920
rect 49973 26911 50031 26917
rect 49973 26877 49985 26911
rect 50019 26908 50031 26911
rect 50338 26908 50344 26920
rect 50019 26880 50344 26908
rect 50019 26877 50031 26880
rect 49973 26871 50031 26877
rect 50338 26868 50344 26880
rect 50396 26868 50402 26920
rect 50706 26868 50712 26920
rect 50764 26908 50770 26920
rect 51442 26908 51448 26920
rect 50764 26880 51448 26908
rect 50764 26868 50770 26880
rect 51442 26868 51448 26880
rect 51500 26908 51506 26920
rect 51629 26911 51687 26917
rect 51629 26908 51641 26911
rect 51500 26880 51641 26908
rect 51500 26868 51506 26880
rect 51629 26877 51641 26880
rect 51675 26877 51687 26911
rect 51629 26871 51687 26877
rect 36596 26812 38976 26840
rect 39669 26843 39727 26849
rect 36596 26800 36602 26812
rect 39669 26809 39681 26843
rect 39715 26840 39727 26843
rect 40034 26840 40040 26852
rect 39715 26812 40040 26840
rect 39715 26809 39727 26812
rect 39669 26803 39727 26809
rect 40034 26800 40040 26812
rect 40092 26840 40098 26852
rect 49234 26840 49240 26852
rect 40092 26812 49240 26840
rect 40092 26800 40098 26812
rect 49234 26800 49240 26812
rect 49292 26840 49298 26852
rect 50154 26840 50160 26852
rect 49292 26812 50160 26840
rect 49292 26800 49298 26812
rect 50154 26800 50160 26812
rect 50212 26800 50218 26852
rect 51074 26800 51080 26852
rect 51132 26840 51138 26852
rect 51132 26812 51177 26840
rect 51132 26800 51138 26812
rect 28644 26744 28994 26772
rect 29273 26775 29331 26781
rect 29273 26741 29285 26775
rect 29319 26772 29331 26775
rect 30650 26772 30656 26784
rect 29319 26744 30656 26772
rect 29319 26741 29331 26744
rect 29273 26735 29331 26741
rect 30650 26732 30656 26744
rect 30708 26732 30714 26784
rect 37369 26775 37427 26781
rect 37369 26741 37381 26775
rect 37415 26772 37427 26775
rect 38746 26772 38752 26784
rect 37415 26744 38752 26772
rect 37415 26741 37427 26744
rect 37369 26735 37427 26741
rect 38746 26732 38752 26744
rect 38804 26732 38810 26784
rect 40129 26775 40187 26781
rect 40129 26741 40141 26775
rect 40175 26772 40187 26775
rect 40402 26772 40408 26784
rect 40175 26744 40408 26772
rect 40175 26741 40187 26744
rect 40129 26735 40187 26741
rect 40402 26732 40408 26744
rect 40460 26732 40466 26784
rect 43717 26775 43775 26781
rect 43717 26741 43729 26775
rect 43763 26772 43775 26775
rect 44082 26772 44088 26784
rect 43763 26744 44088 26772
rect 43763 26741 43775 26744
rect 43717 26735 43775 26741
rect 44082 26732 44088 26744
rect 44140 26732 44146 26784
rect 47670 26732 47676 26784
rect 47728 26772 47734 26784
rect 48133 26775 48191 26781
rect 48133 26772 48145 26775
rect 47728 26744 48145 26772
rect 47728 26732 47734 26744
rect 48133 26741 48145 26744
rect 48179 26772 48191 26775
rect 49326 26772 49332 26784
rect 48179 26744 49332 26772
rect 48179 26741 48191 26744
rect 48133 26735 48191 26741
rect 49326 26732 49332 26744
rect 49384 26732 49390 26784
rect 50338 26732 50344 26784
rect 50396 26772 50402 26784
rect 52454 26772 52460 26784
rect 50396 26744 52460 26772
rect 50396 26732 50402 26744
rect 52454 26732 52460 26744
rect 52512 26732 52518 26784
rect 56962 26732 56968 26784
rect 57020 26772 57026 26784
rect 58069 26775 58127 26781
rect 58069 26772 58081 26775
rect 57020 26744 58081 26772
rect 57020 26732 57026 26744
rect 58069 26741 58081 26744
rect 58115 26741 58127 26775
rect 58069 26735 58127 26741
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 2498 26568 2504 26580
rect 2459 26540 2504 26568
rect 2498 26528 2504 26540
rect 2556 26528 2562 26580
rect 47118 26568 47124 26580
rect 16546 26540 47124 26568
rect 16546 26500 16574 26540
rect 47118 26528 47124 26540
rect 47176 26528 47182 26580
rect 47210 26528 47216 26580
rect 47268 26568 47274 26580
rect 47305 26571 47363 26577
rect 47305 26568 47317 26571
rect 47268 26540 47317 26568
rect 47268 26528 47274 26540
rect 47305 26537 47317 26540
rect 47351 26537 47363 26571
rect 47305 26531 47363 26537
rect 50154 26528 50160 26580
rect 50212 26568 50218 26580
rect 51261 26571 51319 26577
rect 51261 26568 51273 26571
rect 50212 26540 51273 26568
rect 50212 26528 50218 26540
rect 51261 26537 51273 26540
rect 51307 26537 51319 26571
rect 51261 26531 51319 26537
rect 51445 26571 51503 26577
rect 51445 26537 51457 26571
rect 51491 26568 51503 26571
rect 51626 26568 51632 26580
rect 51491 26540 51632 26568
rect 51491 26537 51503 26540
rect 51445 26531 51503 26537
rect 51626 26528 51632 26540
rect 51684 26528 51690 26580
rect 31573 26503 31631 26509
rect 9784 26472 16574 26500
rect 29840 26472 30972 26500
rect 2409 26367 2467 26373
rect 2409 26333 2421 26367
rect 2455 26364 2467 26367
rect 2455 26336 6914 26364
rect 2455 26333 2467 26336
rect 2409 26327 2467 26333
rect 6886 26296 6914 26336
rect 8754 26324 8760 26376
rect 8812 26364 8818 26376
rect 8941 26367 8999 26373
rect 8941 26364 8953 26367
rect 8812 26336 8953 26364
rect 8812 26324 8818 26336
rect 8941 26333 8953 26336
rect 8987 26333 8999 26367
rect 8941 26327 8999 26333
rect 9214 26324 9220 26376
rect 9272 26364 9278 26376
rect 9784 26373 9812 26472
rect 29840 26441 29868 26472
rect 29825 26435 29883 26441
rect 29825 26401 29837 26435
rect 29871 26401 29883 26435
rect 29825 26395 29883 26401
rect 9769 26367 9827 26373
rect 9769 26364 9781 26367
rect 9272 26336 9781 26364
rect 9272 26324 9278 26336
rect 9769 26333 9781 26336
rect 9815 26333 9827 26367
rect 20254 26364 20260 26376
rect 9769 26327 9827 26333
rect 16546 26336 20260 26364
rect 16546 26296 16574 26336
rect 20254 26324 20260 26336
rect 20312 26364 20318 26376
rect 24854 26364 24860 26376
rect 20312 26336 24860 26364
rect 20312 26324 20318 26336
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 29362 26324 29368 26376
rect 29420 26364 29426 26376
rect 29730 26364 29736 26376
rect 29420 26336 29736 26364
rect 29420 26324 29426 26336
rect 29730 26324 29736 26336
rect 29788 26324 29794 26376
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26364 29975 26367
rect 30006 26364 30012 26376
rect 29963 26336 30012 26364
rect 29963 26333 29975 26336
rect 29917 26327 29975 26333
rect 30006 26324 30012 26336
rect 30064 26324 30070 26376
rect 30282 26324 30288 26376
rect 30340 26358 30346 26376
rect 30576 26373 30604 26472
rect 30653 26435 30711 26441
rect 30653 26401 30665 26435
rect 30699 26432 30711 26435
rect 30834 26432 30840 26444
rect 30699 26404 30840 26432
rect 30699 26401 30711 26404
rect 30653 26395 30711 26401
rect 30834 26392 30840 26404
rect 30892 26392 30898 26444
rect 30944 26432 30972 26472
rect 31573 26469 31585 26503
rect 31619 26500 31631 26503
rect 32030 26500 32036 26512
rect 31619 26472 32036 26500
rect 31619 26469 31631 26472
rect 31573 26463 31631 26469
rect 32030 26460 32036 26472
rect 32088 26460 32094 26512
rect 32122 26460 32128 26512
rect 32180 26460 32186 26512
rect 37090 26460 37096 26512
rect 37148 26500 37154 26512
rect 39206 26500 39212 26512
rect 37148 26472 39212 26500
rect 37148 26460 37154 26472
rect 32140 26432 32168 26460
rect 30944 26404 32168 26432
rect 30561 26367 30619 26373
rect 30377 26358 30435 26363
rect 30340 26357 30435 26358
rect 30340 26330 30389 26357
rect 30340 26324 30346 26330
rect 30377 26323 30389 26330
rect 30423 26323 30435 26357
rect 30561 26333 30573 26367
rect 30607 26333 30619 26367
rect 30742 26364 30748 26376
rect 30655 26336 30748 26364
rect 30561 26327 30619 26333
rect 30742 26324 30748 26336
rect 30800 26324 30806 26376
rect 30926 26324 30932 26376
rect 30984 26364 30990 26376
rect 31662 26364 31668 26376
rect 30984 26336 31029 26364
rect 31128 26336 31668 26364
rect 30984 26324 30990 26336
rect 30377 26317 30435 26323
rect 6886 26268 16574 26296
rect 28810 26256 28816 26308
rect 28868 26296 28874 26308
rect 30190 26296 30196 26308
rect 28868 26268 30196 26296
rect 28868 26256 28874 26268
rect 30190 26256 30196 26268
rect 30248 26256 30254 26308
rect 30760 26296 30788 26324
rect 31128 26296 31156 26336
rect 31662 26324 31668 26336
rect 31720 26324 31726 26376
rect 31757 26367 31815 26373
rect 31757 26333 31769 26367
rect 31803 26333 31815 26367
rect 31757 26327 31815 26333
rect 30760 26268 31156 26296
rect 31294 26256 31300 26308
rect 31352 26296 31358 26308
rect 31352 26268 31708 26296
rect 31352 26256 31358 26268
rect 31113 26231 31171 26237
rect 31113 26197 31125 26231
rect 31159 26228 31171 26231
rect 31202 26228 31208 26240
rect 31159 26200 31208 26228
rect 31159 26197 31171 26200
rect 31113 26191 31171 26197
rect 31202 26188 31208 26200
rect 31260 26188 31266 26240
rect 31680 26228 31708 26268
rect 31772 26228 31800 26327
rect 31846 26324 31852 26376
rect 31904 26364 31910 26376
rect 32033 26367 32091 26373
rect 31904 26336 31949 26364
rect 31904 26324 31910 26336
rect 32033 26333 32045 26367
rect 32079 26333 32091 26367
rect 32033 26327 32091 26333
rect 32125 26367 32183 26373
rect 32125 26333 32137 26367
rect 32171 26364 32183 26367
rect 32214 26364 32220 26376
rect 32171 26336 32220 26364
rect 32171 26333 32183 26336
rect 32125 26327 32183 26333
rect 31938 26256 31944 26308
rect 31996 26296 32002 26308
rect 32048 26296 32076 26327
rect 32214 26324 32220 26336
rect 32272 26324 32278 26376
rect 37568 26373 37596 26472
rect 39206 26460 39212 26472
rect 39264 26460 39270 26512
rect 40310 26460 40316 26512
rect 40368 26500 40374 26512
rect 40865 26503 40923 26509
rect 40865 26500 40877 26503
rect 40368 26472 40877 26500
rect 40368 26460 40374 26472
rect 40865 26469 40877 26472
rect 40911 26500 40923 26503
rect 43257 26503 43315 26509
rect 40911 26472 41414 26500
rect 40911 26469 40923 26472
rect 40865 26463 40923 26469
rect 38746 26392 38752 26444
rect 38804 26432 38810 26444
rect 41386 26432 41414 26472
rect 43257 26469 43269 26503
rect 43303 26500 43315 26503
rect 43438 26500 43444 26512
rect 43303 26472 43444 26500
rect 43303 26469 43315 26472
rect 43257 26463 43315 26469
rect 43438 26460 43444 26472
rect 43496 26460 43502 26512
rect 43809 26503 43867 26509
rect 43809 26469 43821 26503
rect 43855 26500 43867 26503
rect 44450 26500 44456 26512
rect 43855 26472 44456 26500
rect 43855 26469 43867 26472
rect 43809 26463 43867 26469
rect 44450 26460 44456 26472
rect 44508 26460 44514 26512
rect 50706 26500 50712 26512
rect 44744 26472 50712 26500
rect 38804 26404 40356 26432
rect 41386 26404 43116 26432
rect 38804 26392 38810 26404
rect 37553 26367 37611 26373
rect 37553 26333 37565 26367
rect 37599 26333 37611 26367
rect 37826 26364 37832 26376
rect 37787 26336 37832 26364
rect 37553 26327 37611 26333
rect 37826 26324 37832 26336
rect 37884 26324 37890 26376
rect 40034 26364 40040 26376
rect 39995 26336 40040 26364
rect 40034 26324 40040 26336
rect 40092 26324 40098 26376
rect 40328 26373 40356 26404
rect 43088 26376 43116 26404
rect 43714 26392 43720 26444
rect 43772 26432 43778 26444
rect 43772 26404 44496 26432
rect 43772 26392 43778 26404
rect 40313 26367 40371 26373
rect 40313 26333 40325 26367
rect 40359 26333 40371 26367
rect 40313 26327 40371 26333
rect 40586 26324 40592 26376
rect 40644 26364 40650 26376
rect 40773 26367 40831 26373
rect 40773 26364 40785 26367
rect 40644 26336 40785 26364
rect 40644 26324 40650 26336
rect 40773 26333 40785 26336
rect 40819 26333 40831 26367
rect 40773 26327 40831 26333
rect 41414 26324 41420 26376
rect 41472 26364 41478 26376
rect 41472 26336 41517 26364
rect 41472 26324 41478 26336
rect 41598 26324 41604 26376
rect 41656 26364 41662 26376
rect 41782 26364 41788 26376
rect 41656 26336 41788 26364
rect 41656 26324 41662 26336
rect 41782 26324 41788 26336
rect 41840 26324 41846 26376
rect 43070 26364 43076 26376
rect 42983 26336 43076 26364
rect 43070 26324 43076 26336
rect 43128 26324 43134 26376
rect 43993 26367 44051 26373
rect 43993 26333 44005 26367
rect 44039 26364 44051 26367
rect 44174 26364 44180 26376
rect 44039 26336 44180 26364
rect 44039 26333 44051 26336
rect 43993 26327 44051 26333
rect 44174 26324 44180 26336
rect 44232 26324 44238 26376
rect 44468 26373 44496 26404
rect 44269 26367 44327 26373
rect 44269 26333 44281 26367
rect 44315 26333 44327 26367
rect 44269 26327 44327 26333
rect 44453 26367 44511 26373
rect 44453 26333 44465 26367
rect 44499 26333 44511 26367
rect 44453 26327 44511 26333
rect 31996 26268 32076 26296
rect 37369 26299 37427 26305
rect 31996 26256 32002 26268
rect 37369 26265 37381 26299
rect 37415 26296 37427 26299
rect 38654 26296 38660 26308
rect 37415 26268 38660 26296
rect 37415 26265 37427 26268
rect 37369 26259 37427 26265
rect 38654 26256 38660 26268
rect 38712 26256 38718 26308
rect 38838 26256 38844 26308
rect 38896 26296 38902 26308
rect 40221 26299 40279 26305
rect 40221 26296 40233 26299
rect 38896 26268 40233 26296
rect 38896 26256 38902 26268
rect 40221 26265 40233 26268
rect 40267 26265 40279 26299
rect 40221 26259 40279 26265
rect 40494 26256 40500 26308
rect 40552 26296 40558 26308
rect 41509 26299 41567 26305
rect 40552 26268 41414 26296
rect 40552 26256 40558 26268
rect 31680 26200 31800 26228
rect 37274 26188 37280 26240
rect 37332 26228 37338 26240
rect 37737 26231 37795 26237
rect 37737 26228 37749 26231
rect 37332 26200 37749 26228
rect 37332 26188 37338 26200
rect 37737 26197 37749 26200
rect 37783 26228 37795 26231
rect 38102 26228 38108 26240
rect 37783 26200 38108 26228
rect 37783 26197 37795 26200
rect 37737 26191 37795 26197
rect 38102 26188 38108 26200
rect 38160 26188 38166 26240
rect 39758 26188 39764 26240
rect 39816 26228 39822 26240
rect 39853 26231 39911 26237
rect 39853 26228 39865 26231
rect 39816 26200 39865 26228
rect 39816 26188 39822 26200
rect 39853 26197 39865 26200
rect 39899 26197 39911 26231
rect 41386 26228 41414 26268
rect 41509 26265 41521 26299
rect 41555 26296 41567 26299
rect 41874 26296 41880 26308
rect 41555 26268 41880 26296
rect 41555 26265 41567 26268
rect 41509 26259 41567 26265
rect 41874 26256 41880 26268
rect 41932 26256 41938 26308
rect 43806 26256 43812 26308
rect 43864 26296 43870 26308
rect 44284 26296 44312 26327
rect 44634 26296 44640 26308
rect 43864 26268 44220 26296
rect 44284 26268 44640 26296
rect 43864 26256 43870 26268
rect 41690 26228 41696 26240
rect 41386 26200 41696 26228
rect 39853 26191 39911 26197
rect 41690 26188 41696 26200
rect 41748 26188 41754 26240
rect 42794 26188 42800 26240
rect 42852 26228 42858 26240
rect 43990 26228 43996 26240
rect 42852 26200 43996 26228
rect 42852 26188 42858 26200
rect 43990 26188 43996 26200
rect 44048 26188 44054 26240
rect 44192 26228 44220 26268
rect 44634 26256 44640 26268
rect 44692 26256 44698 26308
rect 44744 26228 44772 26472
rect 50706 26460 50712 26472
rect 50764 26460 50770 26512
rect 50433 26435 50491 26441
rect 50433 26401 50445 26435
rect 50479 26432 50491 26435
rect 51074 26432 51080 26444
rect 50479 26404 51080 26432
rect 50479 26401 50491 26404
rect 50433 26395 50491 26401
rect 51074 26392 51080 26404
rect 51132 26392 51138 26444
rect 56321 26435 56379 26441
rect 56321 26401 56333 26435
rect 56367 26432 56379 26435
rect 56962 26432 56968 26444
rect 56367 26404 56968 26432
rect 56367 26401 56379 26404
rect 56321 26395 56379 26401
rect 56962 26392 56968 26404
rect 57020 26392 57026 26444
rect 58158 26432 58164 26444
rect 58119 26404 58164 26432
rect 58158 26392 58164 26404
rect 58216 26392 58222 26444
rect 47857 26367 47915 26373
rect 47857 26333 47869 26367
rect 47903 26364 47915 26367
rect 48958 26364 48964 26376
rect 47903 26336 48964 26364
rect 47903 26333 47915 26336
rect 47857 26327 47915 26333
rect 48958 26324 48964 26336
rect 49016 26324 49022 26376
rect 50154 26364 50160 26376
rect 50115 26336 50160 26364
rect 50154 26324 50160 26336
rect 50212 26324 50218 26376
rect 50338 26364 50344 26376
rect 50299 26336 50344 26364
rect 50338 26324 50344 26336
rect 50396 26324 50402 26376
rect 50614 26373 50620 26376
rect 50561 26367 50620 26373
rect 50561 26364 50573 26367
rect 50527 26336 50573 26364
rect 50561 26333 50573 26336
rect 50607 26333 50620 26367
rect 50561 26327 50620 26333
rect 50614 26324 50620 26327
rect 50672 26364 50678 26376
rect 50672 26336 51120 26364
rect 50672 26324 50678 26336
rect 46382 26256 46388 26308
rect 46440 26296 46446 26308
rect 47213 26299 47271 26305
rect 47213 26296 47225 26299
rect 46440 26268 47225 26296
rect 46440 26256 46446 26268
rect 47213 26265 47225 26268
rect 47259 26265 47271 26299
rect 47213 26259 47271 26265
rect 49878 26256 49884 26308
rect 49936 26296 49942 26308
rect 51092 26305 51120 26336
rect 50433 26299 50491 26305
rect 50433 26296 50445 26299
rect 49936 26268 50445 26296
rect 49936 26256 49942 26268
rect 50433 26265 50445 26268
rect 50479 26265 50491 26299
rect 50433 26259 50491 26265
rect 51077 26299 51135 26305
rect 51077 26265 51089 26299
rect 51123 26265 51135 26299
rect 51258 26296 51264 26308
rect 51316 26305 51322 26308
rect 51316 26299 51351 26305
rect 51203 26268 51264 26296
rect 51077 26259 51135 26265
rect 51258 26256 51264 26268
rect 51339 26296 51351 26299
rect 52270 26296 52276 26308
rect 51339 26268 52276 26296
rect 51339 26265 51351 26268
rect 51316 26259 51351 26265
rect 51316 26256 51322 26259
rect 52270 26256 52276 26268
rect 52328 26256 52334 26308
rect 56505 26299 56563 26305
rect 56505 26265 56517 26299
rect 56551 26296 56563 26299
rect 57054 26296 57060 26308
rect 56551 26268 57060 26296
rect 56551 26265 56563 26268
rect 56505 26259 56563 26265
rect 57054 26256 57060 26268
rect 57112 26256 57118 26308
rect 44192 26200 44772 26228
rect 47670 26188 47676 26240
rect 47728 26228 47734 26240
rect 47949 26231 48007 26237
rect 47949 26228 47961 26231
rect 47728 26200 47961 26228
rect 47728 26188 47734 26200
rect 47949 26197 47961 26200
rect 47995 26228 48007 26231
rect 48038 26228 48044 26240
rect 47995 26200 48044 26228
rect 47995 26197 48007 26200
rect 47949 26191 48007 26197
rect 48038 26188 48044 26200
rect 48096 26188 48102 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 37366 25984 37372 26036
rect 37424 26024 37430 26036
rect 40862 26024 40868 26036
rect 37424 25996 40868 26024
rect 37424 25984 37430 25996
rect 40862 25984 40868 25996
rect 40920 25984 40926 26036
rect 41417 26027 41475 26033
rect 41417 25993 41429 26027
rect 41463 26024 41475 26027
rect 43714 26024 43720 26036
rect 41463 25996 43720 26024
rect 41463 25993 41475 25996
rect 41417 25987 41475 25993
rect 43714 25984 43720 25996
rect 43772 25984 43778 26036
rect 44729 26027 44787 26033
rect 44729 25993 44741 26027
rect 44775 26024 44787 26027
rect 46290 26024 46296 26036
rect 44775 25996 46296 26024
rect 44775 25993 44787 25996
rect 44729 25987 44787 25993
rect 46290 25984 46296 25996
rect 46348 25984 46354 26036
rect 49234 25984 49240 26036
rect 49292 26024 49298 26036
rect 51258 26024 51264 26036
rect 49292 25996 51264 26024
rect 49292 25984 49298 25996
rect 51258 25984 51264 25996
rect 51316 25984 51322 26036
rect 57054 26024 57060 26036
rect 57015 25996 57060 26024
rect 57054 25984 57060 25996
rect 57112 25984 57118 26036
rect 2682 25916 2688 25968
rect 2740 25956 2746 25968
rect 7745 25959 7803 25965
rect 7745 25956 7757 25959
rect 2740 25928 7757 25956
rect 2740 25916 2746 25928
rect 7745 25925 7757 25928
rect 7791 25925 7803 25959
rect 7745 25919 7803 25925
rect 9858 25916 9864 25968
rect 9916 25956 9922 25968
rect 16574 25956 16580 25968
rect 9916 25928 16580 25956
rect 9916 25916 9922 25928
rect 16574 25916 16580 25928
rect 16632 25956 16638 25968
rect 39574 25956 39580 25968
rect 16632 25928 39580 25956
rect 16632 25916 16638 25928
rect 39574 25916 39580 25928
rect 39632 25916 39638 25968
rect 39684 25919 39804 25922
rect 39684 25913 39819 25919
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25888 8171 25891
rect 8754 25888 8760 25900
rect 8159 25860 8760 25888
rect 8159 25857 8171 25860
rect 8113 25851 8171 25857
rect 8754 25848 8760 25860
rect 8812 25848 8818 25900
rect 30374 25888 30380 25900
rect 30335 25860 30380 25888
rect 30374 25848 30380 25860
rect 30432 25848 30438 25900
rect 30469 25891 30527 25897
rect 30469 25857 30481 25891
rect 30515 25857 30527 25891
rect 30650 25888 30656 25900
rect 30611 25860 30656 25888
rect 30469 25851 30527 25857
rect 9490 25780 9496 25832
rect 9548 25820 9554 25832
rect 9585 25823 9643 25829
rect 9585 25820 9597 25823
rect 9548 25792 9597 25820
rect 9548 25780 9554 25792
rect 9585 25789 9597 25792
rect 9631 25820 9643 25823
rect 26970 25820 26976 25832
rect 9631 25792 26976 25820
rect 9631 25789 9643 25792
rect 9585 25783 9643 25789
rect 26970 25780 26976 25792
rect 27028 25780 27034 25832
rect 29546 25780 29552 25832
rect 29604 25820 29610 25832
rect 30484 25820 30512 25851
rect 30650 25848 30656 25860
rect 30708 25848 30714 25900
rect 30745 25891 30803 25897
rect 30745 25857 30757 25891
rect 30791 25857 30803 25891
rect 31202 25888 31208 25900
rect 31163 25860 31208 25888
rect 30745 25851 30803 25857
rect 29604 25792 30512 25820
rect 30760 25820 30788 25851
rect 31202 25848 31208 25860
rect 31260 25848 31266 25900
rect 31389 25891 31447 25897
rect 31389 25857 31401 25891
rect 31435 25888 31447 25891
rect 31478 25888 31484 25900
rect 31435 25860 31484 25888
rect 31435 25857 31447 25860
rect 31389 25851 31447 25857
rect 31478 25848 31484 25860
rect 31536 25848 31542 25900
rect 37274 25888 37280 25900
rect 37235 25860 37280 25888
rect 37274 25848 37280 25860
rect 37332 25848 37338 25900
rect 37550 25888 37556 25900
rect 37511 25860 37556 25888
rect 37550 25848 37556 25860
rect 37608 25848 37614 25900
rect 37642 25848 37648 25900
rect 37700 25888 37706 25900
rect 37737 25891 37795 25897
rect 37737 25888 37749 25891
rect 37700 25860 37749 25888
rect 37700 25848 37706 25860
rect 37737 25857 37749 25860
rect 37783 25857 37795 25891
rect 38010 25888 38016 25900
rect 37971 25860 38016 25888
rect 37737 25851 37795 25857
rect 38010 25848 38016 25860
rect 38068 25848 38074 25900
rect 38930 25888 38936 25900
rect 38891 25860 38936 25888
rect 38930 25848 38936 25860
rect 38988 25848 38994 25900
rect 39482 25848 39488 25900
rect 39540 25888 39546 25900
rect 39684 25894 39773 25913
rect 39684 25888 39712 25894
rect 39540 25860 39712 25888
rect 39761 25879 39773 25894
rect 39807 25879 39819 25913
rect 39850 25882 39856 25934
rect 39908 25922 39914 25934
rect 39908 25894 39953 25922
rect 40310 25916 40316 25968
rect 40368 25956 40374 25968
rect 40368 25928 51074 25956
rect 40368 25916 40374 25928
rect 40034 25897 40040 25900
rect 39908 25882 39914 25894
rect 39991 25891 40040 25897
rect 39761 25873 39819 25879
rect 39540 25848 39546 25860
rect 39991 25857 40003 25891
rect 40037 25857 40040 25891
rect 39991 25851 40040 25857
rect 40034 25848 40040 25851
rect 40092 25848 40098 25900
rect 40129 25891 40187 25897
rect 40129 25857 40141 25891
rect 40175 25857 40187 25891
rect 40129 25851 40187 25857
rect 40221 25891 40279 25897
rect 40221 25857 40233 25891
rect 40267 25888 40279 25891
rect 40586 25888 40592 25900
rect 40267 25860 40592 25888
rect 40267 25857 40279 25860
rect 40221 25851 40279 25857
rect 32858 25820 32864 25832
rect 30760 25792 32864 25820
rect 29604 25780 29610 25792
rect 32858 25780 32864 25792
rect 32916 25780 32922 25832
rect 38746 25820 38752 25832
rect 38707 25792 38752 25820
rect 38746 25780 38752 25792
rect 38804 25780 38810 25832
rect 38838 25780 38844 25832
rect 38896 25820 38902 25832
rect 39025 25823 39083 25829
rect 38896 25792 38941 25820
rect 38896 25780 38902 25792
rect 39025 25789 39037 25823
rect 39071 25789 39083 25823
rect 40144 25820 40172 25851
rect 40586 25848 40592 25860
rect 40644 25848 40650 25900
rect 40773 25891 40831 25897
rect 40773 25857 40785 25891
rect 40819 25888 40831 25891
rect 40862 25888 40868 25900
rect 40819 25860 40868 25888
rect 40819 25857 40831 25860
rect 40773 25851 40831 25857
rect 40862 25848 40868 25860
rect 40920 25848 40926 25900
rect 41598 25888 41604 25900
rect 41559 25860 41604 25888
rect 41598 25848 41604 25860
rect 41656 25848 41662 25900
rect 41782 25888 41788 25900
rect 41743 25860 41788 25888
rect 41782 25848 41788 25860
rect 41840 25848 41846 25900
rect 41877 25891 41935 25897
rect 41877 25857 41889 25891
rect 41923 25857 41935 25891
rect 43438 25888 43444 25900
rect 43399 25860 43444 25888
rect 41877 25851 41935 25857
rect 40310 25820 40316 25832
rect 40144 25792 40316 25820
rect 39025 25783 39083 25789
rect 37829 25755 37887 25761
rect 37829 25721 37841 25755
rect 37875 25752 37887 25755
rect 38856 25752 38884 25780
rect 37875 25724 38884 25752
rect 37875 25721 37887 25724
rect 37829 25715 37887 25721
rect 29362 25644 29368 25696
rect 29420 25684 29426 25696
rect 30193 25687 30251 25693
rect 30193 25684 30205 25687
rect 29420 25656 30205 25684
rect 29420 25644 29426 25656
rect 30193 25653 30205 25656
rect 30239 25653 30251 25687
rect 30193 25647 30251 25653
rect 31018 25644 31024 25696
rect 31076 25684 31082 25696
rect 31205 25687 31263 25693
rect 31205 25684 31217 25687
rect 31076 25656 31217 25684
rect 31076 25644 31082 25656
rect 31205 25653 31217 25656
rect 31251 25653 31263 25687
rect 31205 25647 31263 25653
rect 38286 25644 38292 25696
rect 38344 25684 38350 25696
rect 38565 25687 38623 25693
rect 38565 25684 38577 25687
rect 38344 25656 38577 25684
rect 38344 25644 38350 25656
rect 38565 25653 38577 25656
rect 38611 25653 38623 25687
rect 39040 25684 39068 25783
rect 40310 25780 40316 25792
rect 40368 25780 40374 25832
rect 41414 25820 41420 25832
rect 41386 25780 41420 25820
rect 41472 25820 41478 25832
rect 41892 25820 41920 25851
rect 43438 25848 43444 25860
rect 43496 25848 43502 25900
rect 43530 25848 43536 25900
rect 43588 25888 43594 25900
rect 43625 25891 43683 25897
rect 43625 25888 43637 25891
rect 43588 25860 43637 25888
rect 43588 25848 43594 25860
rect 43625 25857 43637 25860
rect 43671 25857 43683 25891
rect 43625 25851 43683 25857
rect 43809 25891 43867 25897
rect 43809 25857 43821 25891
rect 43855 25888 43867 25891
rect 44358 25888 44364 25900
rect 43855 25860 44364 25888
rect 43855 25857 43867 25860
rect 43809 25851 43867 25857
rect 44358 25848 44364 25860
rect 44416 25888 44422 25900
rect 44453 25891 44511 25897
rect 44453 25888 44465 25891
rect 44416 25860 44465 25888
rect 44416 25848 44422 25860
rect 44453 25857 44465 25860
rect 44499 25857 44511 25891
rect 48866 25888 48872 25900
rect 48827 25860 48872 25888
rect 44453 25851 44511 25857
rect 48866 25848 48872 25860
rect 48924 25848 48930 25900
rect 49053 25891 49111 25897
rect 49053 25857 49065 25891
rect 49099 25888 49111 25891
rect 49694 25888 49700 25900
rect 49099 25860 49700 25888
rect 49099 25857 49111 25860
rect 49053 25851 49111 25857
rect 44266 25820 44272 25832
rect 41472 25792 41920 25820
rect 44227 25792 44272 25820
rect 41472 25780 41478 25792
rect 44266 25780 44272 25792
rect 44324 25780 44330 25832
rect 44821 25823 44879 25829
rect 44821 25820 44833 25823
rect 44376 25792 44833 25820
rect 39577 25755 39635 25761
rect 39577 25721 39589 25755
rect 39623 25752 39635 25755
rect 41386 25752 41414 25780
rect 39623 25724 41414 25752
rect 39623 25721 39635 25724
rect 39577 25715 39635 25721
rect 44082 25712 44088 25764
rect 44140 25752 44146 25764
rect 44376 25752 44404 25792
rect 44821 25789 44833 25792
rect 44867 25789 44879 25823
rect 49068 25820 49096 25851
rect 49694 25848 49700 25860
rect 49752 25848 49758 25900
rect 51046 25888 51074 25928
rect 56321 25891 56379 25897
rect 56321 25888 56333 25891
rect 51046 25860 56333 25888
rect 56321 25857 56333 25860
rect 56367 25857 56379 25891
rect 56321 25851 56379 25857
rect 56965 25891 57023 25897
rect 56965 25857 56977 25891
rect 57011 25888 57023 25891
rect 57422 25888 57428 25900
rect 57011 25860 57428 25888
rect 57011 25857 57023 25860
rect 56965 25851 57023 25857
rect 57422 25848 57428 25860
rect 57480 25848 57486 25900
rect 44821 25783 44879 25789
rect 47780 25792 49096 25820
rect 44140 25724 44404 25752
rect 44140 25712 44146 25724
rect 47780 25696 47808 25792
rect 40402 25684 40408 25696
rect 39040 25656 40408 25684
rect 38565 25647 38623 25653
rect 40402 25644 40408 25656
rect 40460 25644 40466 25696
rect 40678 25644 40684 25696
rect 40736 25684 40742 25696
rect 40865 25687 40923 25693
rect 40865 25684 40877 25687
rect 40736 25656 40877 25684
rect 40736 25644 40742 25656
rect 40865 25653 40877 25656
rect 40911 25653 40923 25687
rect 40865 25647 40923 25653
rect 41690 25644 41696 25696
rect 41748 25684 41754 25696
rect 47762 25684 47768 25696
rect 41748 25656 47768 25684
rect 41748 25644 41754 25656
rect 47762 25644 47768 25656
rect 47820 25644 47826 25696
rect 49234 25684 49240 25696
rect 49195 25656 49240 25684
rect 49234 25644 49240 25656
rect 49292 25644 49298 25696
rect 56413 25687 56471 25693
rect 56413 25653 56425 25687
rect 56459 25684 56471 25687
rect 56502 25684 56508 25696
rect 56459 25656 56508 25684
rect 56459 25653 56471 25656
rect 56413 25647 56471 25653
rect 56502 25644 56508 25656
rect 56560 25644 56566 25696
rect 58066 25684 58072 25696
rect 58027 25656 58072 25684
rect 58066 25644 58072 25656
rect 58124 25644 58130 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 39301 25483 39359 25489
rect 39301 25449 39313 25483
rect 39347 25480 39359 25483
rect 40034 25480 40040 25492
rect 39347 25452 40040 25480
rect 39347 25449 39359 25452
rect 39301 25443 39359 25449
rect 40034 25440 40040 25452
rect 40092 25440 40098 25492
rect 42794 25440 42800 25492
rect 42852 25440 42858 25492
rect 44269 25483 44327 25489
rect 44269 25449 44281 25483
rect 44315 25480 44327 25483
rect 44358 25480 44364 25492
rect 44315 25452 44364 25480
rect 44315 25449 44327 25452
rect 44269 25443 44327 25449
rect 44358 25440 44364 25452
rect 44416 25480 44422 25492
rect 45278 25480 45284 25492
rect 44416 25452 45284 25480
rect 44416 25440 44422 25452
rect 45278 25440 45284 25452
rect 45336 25440 45342 25492
rect 36817 25415 36875 25421
rect 36817 25381 36829 25415
rect 36863 25412 36875 25415
rect 36863 25384 37412 25412
rect 36863 25381 36875 25384
rect 36817 25375 36875 25381
rect 36541 25347 36599 25353
rect 36541 25313 36553 25347
rect 36587 25344 36599 25347
rect 37090 25344 37096 25356
rect 36587 25316 37096 25344
rect 36587 25313 36599 25316
rect 36541 25307 36599 25313
rect 37090 25304 37096 25316
rect 37148 25304 37154 25356
rect 37384 25353 37412 25384
rect 38746 25372 38752 25424
rect 38804 25412 38810 25424
rect 39114 25412 39120 25424
rect 38804 25384 39120 25412
rect 38804 25372 38810 25384
rect 39114 25372 39120 25384
rect 39172 25372 39178 25424
rect 40126 25372 40132 25424
rect 40184 25412 40190 25424
rect 40957 25415 41015 25421
rect 40184 25384 40264 25412
rect 40184 25372 40190 25384
rect 37369 25347 37427 25353
rect 37369 25313 37381 25347
rect 37415 25313 37427 25347
rect 39482 25344 39488 25356
rect 37369 25307 37427 25313
rect 38304 25316 39488 25344
rect 38304 25288 38332 25316
rect 39482 25304 39488 25316
rect 39540 25344 39546 25356
rect 40236 25353 40264 25384
rect 40957 25381 40969 25415
rect 41003 25381 41015 25415
rect 40957 25375 41015 25381
rect 40037 25347 40095 25353
rect 40037 25344 40049 25347
rect 39540 25316 40049 25344
rect 39540 25304 39546 25316
rect 40037 25313 40049 25316
rect 40083 25313 40095 25347
rect 40037 25307 40095 25313
rect 40212 25347 40270 25353
rect 40212 25313 40224 25347
rect 40258 25344 40270 25347
rect 40972 25344 41000 25375
rect 40258 25316 41000 25344
rect 40258 25313 40270 25316
rect 40212 25307 40270 25313
rect 8754 25236 8760 25288
rect 8812 25276 8818 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8812 25248 8953 25276
rect 8812 25236 8818 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 36449 25279 36507 25285
rect 36449 25245 36461 25279
rect 36495 25276 36507 25279
rect 37274 25276 37280 25288
rect 36495 25248 37280 25276
rect 36495 25245 36507 25248
rect 36449 25239 36507 25245
rect 37274 25236 37280 25248
rect 37332 25236 37338 25288
rect 37461 25279 37519 25285
rect 37461 25245 37473 25279
rect 37507 25276 37519 25279
rect 38010 25276 38016 25288
rect 37507 25248 38016 25276
rect 37507 25245 37519 25248
rect 37461 25239 37519 25245
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 38473 25279 38531 25285
rect 38473 25245 38485 25279
rect 38519 25245 38531 25279
rect 38473 25239 38531 25245
rect 9858 25208 9864 25220
rect 9819 25180 9864 25208
rect 9858 25168 9864 25180
rect 9916 25168 9922 25220
rect 38488 25208 38516 25239
rect 38838 25236 38844 25288
rect 38896 25276 38902 25288
rect 38933 25279 38991 25285
rect 38933 25276 38945 25279
rect 38896 25248 38945 25276
rect 38896 25236 38902 25248
rect 38933 25245 38945 25248
rect 38979 25245 38991 25279
rect 39114 25276 39120 25288
rect 39075 25248 39120 25276
rect 38933 25239 38991 25245
rect 39114 25236 39120 25248
rect 39172 25236 39178 25288
rect 40129 25279 40187 25285
rect 40129 25278 40141 25279
rect 40052 25250 40141 25278
rect 39758 25208 39764 25220
rect 38488 25180 39764 25208
rect 39758 25168 39764 25180
rect 39816 25208 39822 25220
rect 40052 25208 40080 25250
rect 40129 25245 40141 25250
rect 40175 25245 40187 25279
rect 40310 25276 40316 25288
rect 40271 25248 40316 25276
rect 40129 25239 40187 25245
rect 40310 25236 40316 25248
rect 40368 25236 40374 25288
rect 40494 25236 40500 25288
rect 40552 25276 40558 25288
rect 41138 25276 41144 25288
rect 40552 25248 41144 25276
rect 40552 25236 40558 25248
rect 41138 25236 41144 25248
rect 41196 25236 41202 25288
rect 41230 25236 41236 25288
rect 41288 25276 41294 25288
rect 41785 25279 41843 25285
rect 41785 25276 41797 25279
rect 41288 25248 41797 25276
rect 41288 25236 41294 25248
rect 41785 25245 41797 25248
rect 41831 25245 41843 25279
rect 42702 25276 42708 25288
rect 42663 25248 42708 25276
rect 41785 25239 41843 25245
rect 42702 25236 42708 25248
rect 42760 25236 42766 25288
rect 42812 25285 42840 25440
rect 44174 25372 44180 25424
rect 44232 25412 44238 25424
rect 44453 25415 44511 25421
rect 44453 25412 44465 25415
rect 44232 25384 44465 25412
rect 44232 25372 44238 25384
rect 44453 25381 44465 25384
rect 44499 25381 44511 25415
rect 58066 25412 58072 25424
rect 44453 25375 44511 25381
rect 56336 25384 58072 25412
rect 47670 25344 47676 25356
rect 47136 25316 47676 25344
rect 42797 25279 42855 25285
rect 42797 25245 42809 25279
rect 42843 25245 42855 25279
rect 42797 25239 42855 25245
rect 42886 25236 42892 25288
rect 42944 25276 42950 25288
rect 42944 25248 42989 25276
rect 42944 25236 42950 25248
rect 43070 25236 43076 25288
rect 43128 25276 43134 25288
rect 43128 25248 43173 25276
rect 43128 25236 43134 25248
rect 43438 25236 43444 25288
rect 43496 25276 43502 25288
rect 47136 25285 47164 25316
rect 47670 25304 47676 25316
rect 47728 25304 47734 25356
rect 56336 25353 56364 25384
rect 58066 25372 58072 25384
rect 58124 25372 58130 25424
rect 56321 25347 56379 25353
rect 56321 25313 56333 25347
rect 56367 25313 56379 25347
rect 56502 25344 56508 25356
rect 56463 25316 56508 25344
rect 56321 25307 56379 25313
rect 56502 25304 56508 25316
rect 56560 25304 56566 25356
rect 58158 25344 58164 25356
rect 58119 25316 58164 25344
rect 58158 25304 58164 25316
rect 58216 25304 58222 25356
rect 45005 25279 45063 25285
rect 45005 25276 45017 25279
rect 43496 25248 45017 25276
rect 43496 25236 43502 25248
rect 45005 25245 45017 25248
rect 45051 25245 45063 25279
rect 45005 25239 45063 25245
rect 47121 25279 47179 25285
rect 47121 25245 47133 25279
rect 47167 25245 47179 25279
rect 47121 25239 47179 25245
rect 47305 25279 47363 25285
rect 47305 25245 47317 25279
rect 47351 25245 47363 25279
rect 47762 25276 47768 25288
rect 47723 25248 47768 25276
rect 47305 25239 47363 25245
rect 39816 25180 40080 25208
rect 40865 25211 40923 25217
rect 39816 25168 39822 25180
rect 40865 25177 40877 25211
rect 40911 25177 40923 25211
rect 40865 25171 40923 25177
rect 37826 25140 37832 25152
rect 37787 25112 37832 25140
rect 37826 25100 37832 25112
rect 37884 25100 37890 25152
rect 38473 25143 38531 25149
rect 38473 25109 38485 25143
rect 38519 25140 38531 25143
rect 39114 25140 39120 25152
rect 38519 25112 39120 25140
rect 38519 25109 38531 25112
rect 38473 25103 38531 25109
rect 39114 25100 39120 25112
rect 39172 25100 39178 25152
rect 39853 25143 39911 25149
rect 39853 25109 39865 25143
rect 39899 25140 39911 25143
rect 40218 25140 40224 25152
rect 39899 25112 40224 25140
rect 39899 25109 39911 25112
rect 39853 25103 39911 25109
rect 40218 25100 40224 25112
rect 40276 25100 40282 25152
rect 40880 25140 40908 25171
rect 40954 25168 40960 25220
rect 41012 25208 41018 25220
rect 41049 25211 41107 25217
rect 41049 25208 41061 25211
rect 41012 25180 41061 25208
rect 41012 25168 41018 25180
rect 41049 25177 41061 25180
rect 41095 25177 41107 25211
rect 41966 25208 41972 25220
rect 41927 25180 41972 25208
rect 41049 25171 41107 25177
rect 41966 25168 41972 25180
rect 42024 25168 42030 25220
rect 44082 25208 44088 25220
rect 44043 25180 44088 25208
rect 44082 25168 44088 25180
rect 44140 25168 44146 25220
rect 47320 25208 47348 25239
rect 47762 25236 47768 25248
rect 47820 25236 47826 25288
rect 47949 25279 48007 25285
rect 47949 25245 47961 25279
rect 47995 25276 48007 25279
rect 48866 25276 48872 25288
rect 47995 25248 48872 25276
rect 47995 25245 48007 25248
rect 47949 25239 48007 25245
rect 47964 25208 47992 25239
rect 48866 25236 48872 25248
rect 48924 25236 48930 25288
rect 47320 25180 47992 25208
rect 41414 25140 41420 25152
rect 40880 25112 41420 25140
rect 41414 25100 41420 25112
rect 41472 25100 41478 25152
rect 41782 25100 41788 25152
rect 41840 25140 41846 25152
rect 41984 25140 42012 25168
rect 41840 25112 42012 25140
rect 42429 25143 42487 25149
rect 41840 25100 41846 25112
rect 42429 25109 42441 25143
rect 42475 25140 42487 25143
rect 43990 25140 43996 25152
rect 42475 25112 43996 25140
rect 42475 25109 42487 25112
rect 42429 25103 42487 25109
rect 43990 25100 43996 25112
rect 44048 25100 44054 25152
rect 44266 25100 44272 25152
rect 44324 25149 44330 25152
rect 44324 25143 44343 25149
rect 44331 25109 44343 25143
rect 45186 25140 45192 25152
rect 45147 25112 45192 25140
rect 44324 25103 44343 25109
rect 44324 25100 44330 25103
rect 45186 25100 45192 25112
rect 45244 25100 45250 25152
rect 47302 25140 47308 25152
rect 47263 25112 47308 25140
rect 47302 25100 47308 25112
rect 47360 25100 47366 25152
rect 47670 25100 47676 25152
rect 47728 25140 47734 25152
rect 47857 25143 47915 25149
rect 47857 25140 47869 25143
rect 47728 25112 47869 25140
rect 47728 25100 47734 25112
rect 47857 25109 47869 25112
rect 47903 25109 47915 25143
rect 47857 25103 47915 25109
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 38654 24896 38660 24948
rect 38712 24936 38718 24948
rect 38712 24908 38757 24936
rect 38712 24896 38718 24908
rect 38838 24896 38844 24948
rect 38896 24936 38902 24948
rect 39419 24939 39477 24945
rect 39419 24936 39431 24939
rect 38896 24908 39431 24936
rect 38896 24896 38902 24908
rect 39419 24905 39431 24908
rect 39465 24936 39477 24939
rect 41414 24936 41420 24948
rect 39465 24908 41420 24936
rect 39465 24905 39477 24908
rect 39419 24899 39477 24905
rect 41414 24896 41420 24908
rect 41472 24896 41478 24948
rect 42886 24936 42892 24948
rect 42812 24908 42892 24936
rect 37369 24871 37427 24877
rect 37369 24837 37381 24871
rect 37415 24868 37427 24871
rect 37826 24868 37832 24880
rect 37415 24840 37832 24868
rect 37415 24837 37427 24840
rect 37369 24831 37427 24837
rect 37826 24828 37832 24840
rect 37884 24828 37890 24880
rect 39209 24871 39267 24877
rect 39209 24868 39221 24871
rect 38488 24840 39221 24868
rect 2314 24800 2320 24812
rect 2275 24772 2320 24800
rect 2314 24760 2320 24772
rect 2372 24800 2378 24812
rect 8570 24800 8576 24812
rect 2372 24772 8576 24800
rect 2372 24760 2378 24772
rect 8570 24760 8576 24772
rect 8628 24760 8634 24812
rect 8754 24800 8760 24812
rect 8715 24772 8760 24800
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 37550 24800 37556 24812
rect 37511 24772 37556 24800
rect 37550 24760 37556 24772
rect 37608 24760 37614 24812
rect 37645 24803 37703 24809
rect 37645 24769 37657 24803
rect 37691 24800 37703 24803
rect 38102 24800 38108 24812
rect 37691 24772 38108 24800
rect 37691 24769 37703 24772
rect 37645 24763 37703 24769
rect 38102 24760 38108 24772
rect 38160 24760 38166 24812
rect 38488 24809 38516 24840
rect 39209 24837 39221 24840
rect 39255 24868 39267 24871
rect 40494 24868 40500 24880
rect 39255 24840 40500 24868
rect 39255 24837 39267 24840
rect 39209 24831 39267 24837
rect 40494 24828 40500 24840
rect 40552 24828 40558 24880
rect 41230 24868 41236 24880
rect 41191 24840 41236 24868
rect 41230 24828 41236 24840
rect 41288 24828 41294 24880
rect 38473 24803 38531 24809
rect 38473 24769 38485 24803
rect 38519 24769 38531 24803
rect 38749 24803 38807 24809
rect 38749 24800 38761 24803
rect 38473 24763 38531 24769
rect 38626 24772 38761 24800
rect 9030 24732 9036 24744
rect 8991 24704 9036 24732
rect 9030 24692 9036 24704
rect 9088 24692 9094 24744
rect 38626 24732 38654 24772
rect 38749 24769 38761 24772
rect 38795 24800 38807 24803
rect 38838 24800 38844 24812
rect 38795 24772 38844 24800
rect 38795 24769 38807 24772
rect 38749 24763 38807 24769
rect 38838 24760 38844 24772
rect 38896 24760 38902 24812
rect 39114 24760 39120 24812
rect 39172 24800 39178 24812
rect 40221 24803 40279 24809
rect 40221 24800 40233 24803
rect 39172 24772 40233 24800
rect 39172 24760 39178 24772
rect 40221 24769 40233 24772
rect 40267 24769 40279 24803
rect 41046 24800 41052 24812
rect 41007 24772 41052 24800
rect 40221 24763 40279 24769
rect 41046 24760 41052 24772
rect 41104 24760 41110 24812
rect 41325 24803 41383 24809
rect 41325 24769 41337 24803
rect 41371 24769 41383 24803
rect 41325 24763 41383 24769
rect 40310 24732 40316 24744
rect 37660 24704 38654 24732
rect 40271 24704 40316 24732
rect 37660 24673 37688 24704
rect 40310 24692 40316 24704
rect 40368 24692 40374 24744
rect 37645 24667 37703 24673
rect 37645 24633 37657 24667
rect 37691 24633 37703 24667
rect 37645 24627 37703 24633
rect 38654 24624 38660 24676
rect 38712 24664 38718 24676
rect 40954 24664 40960 24676
rect 38712 24636 40960 24664
rect 38712 24624 38718 24636
rect 1857 24599 1915 24605
rect 1857 24565 1869 24599
rect 1903 24596 1915 24599
rect 1946 24596 1952 24608
rect 1903 24568 1952 24596
rect 1903 24565 1915 24568
rect 1857 24559 1915 24565
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 2130 24556 2136 24608
rect 2188 24596 2194 24608
rect 2409 24599 2467 24605
rect 2409 24596 2421 24599
rect 2188 24568 2421 24596
rect 2188 24556 2194 24568
rect 2409 24565 2421 24568
rect 2455 24565 2467 24599
rect 2409 24559 2467 24565
rect 38473 24599 38531 24605
rect 38473 24565 38485 24599
rect 38519 24596 38531 24599
rect 39298 24596 39304 24608
rect 38519 24568 39304 24596
rect 38519 24565 38531 24568
rect 38473 24559 38531 24565
rect 39298 24556 39304 24568
rect 39356 24556 39362 24608
rect 39408 24605 39436 24636
rect 40954 24624 40960 24636
rect 41012 24664 41018 24676
rect 41340 24664 41368 24763
rect 41414 24760 41420 24812
rect 41472 24800 41478 24812
rect 42613 24803 42671 24809
rect 42613 24800 42625 24803
rect 41472 24772 41517 24800
rect 41616 24772 42625 24800
rect 41472 24760 41478 24772
rect 41616 24673 41644 24772
rect 42613 24769 42625 24772
rect 42659 24800 42671 24803
rect 42812 24800 42840 24908
rect 42886 24896 42892 24908
rect 42944 24896 42950 24948
rect 44453 24939 44511 24945
rect 44453 24905 44465 24939
rect 44499 24936 44511 24939
rect 45186 24936 45192 24948
rect 44499 24908 45192 24936
rect 44499 24905 44511 24908
rect 44453 24899 44511 24905
rect 45186 24896 45192 24908
rect 45244 24896 45250 24948
rect 47210 24896 47216 24948
rect 47268 24936 47274 24948
rect 47949 24939 48007 24945
rect 47949 24936 47961 24939
rect 47268 24908 47961 24936
rect 47268 24896 47274 24908
rect 47949 24905 47961 24908
rect 47995 24905 48007 24939
rect 47949 24899 48007 24905
rect 44634 24828 44640 24880
rect 44692 24868 44698 24880
rect 46290 24868 46296 24880
rect 44692 24840 46296 24868
rect 44692 24828 44698 24840
rect 46290 24828 46296 24840
rect 46348 24828 46354 24880
rect 42659 24772 42840 24800
rect 42889 24803 42947 24809
rect 42659 24769 42671 24772
rect 42613 24763 42671 24769
rect 42889 24769 42901 24803
rect 42935 24800 42947 24803
rect 42978 24800 42984 24812
rect 42935 24772 42984 24800
rect 42935 24769 42947 24772
rect 42889 24763 42947 24769
rect 42978 24760 42984 24772
rect 43036 24760 43042 24812
rect 43441 24803 43499 24809
rect 43441 24769 43453 24803
rect 43487 24769 43499 24803
rect 43441 24763 43499 24769
rect 41874 24692 41880 24744
rect 41932 24732 41938 24744
rect 43456 24732 43484 24763
rect 44542 24732 44548 24744
rect 41932 24704 43484 24732
rect 44503 24704 44548 24732
rect 41932 24692 41938 24704
rect 44542 24692 44548 24704
rect 44600 24692 44606 24744
rect 44652 24741 44680 24828
rect 45278 24800 45284 24812
rect 45239 24772 45284 24800
rect 45278 24760 45284 24772
rect 45336 24760 45342 24812
rect 46382 24760 46388 24812
rect 46440 24800 46446 24812
rect 46496 24803 46554 24809
rect 46496 24800 46508 24803
rect 46440 24772 46508 24800
rect 46440 24760 46446 24772
rect 46496 24769 46508 24772
rect 46542 24769 46554 24803
rect 46661 24803 46719 24809
rect 46661 24800 46673 24803
rect 46496 24763 46554 24769
rect 46584 24772 46673 24800
rect 44637 24735 44695 24741
rect 44637 24701 44649 24735
rect 44683 24701 44695 24735
rect 44637 24695 44695 24701
rect 41012 24636 41368 24664
rect 41601 24667 41659 24673
rect 41012 24624 41018 24636
rect 41601 24633 41613 24667
rect 41647 24633 41659 24667
rect 42794 24664 42800 24676
rect 41601 24627 41659 24633
rect 42352 24636 42800 24664
rect 39393 24599 39451 24605
rect 39393 24565 39405 24599
rect 39439 24565 39451 24599
rect 39393 24559 39451 24565
rect 39577 24599 39635 24605
rect 39577 24565 39589 24599
rect 39623 24596 39635 24599
rect 40126 24596 40132 24608
rect 39623 24568 40132 24596
rect 39623 24565 39635 24568
rect 39577 24559 39635 24565
rect 40126 24556 40132 24568
rect 40184 24556 40190 24608
rect 40497 24599 40555 24605
rect 40497 24565 40509 24599
rect 40543 24596 40555 24599
rect 42352 24596 42380 24636
rect 42794 24624 42800 24636
rect 42852 24624 42858 24676
rect 43622 24664 43628 24676
rect 43583 24636 43628 24664
rect 43622 24624 43628 24636
rect 43680 24624 43686 24676
rect 43990 24624 43996 24676
rect 44048 24664 44054 24676
rect 44726 24664 44732 24676
rect 44048 24636 44732 24664
rect 44048 24624 44054 24636
rect 44726 24624 44732 24636
rect 44784 24664 44790 24676
rect 44784 24636 45416 24664
rect 44784 24624 44790 24636
rect 40543 24568 42380 24596
rect 42429 24599 42487 24605
rect 40543 24565 40555 24568
rect 40497 24559 40555 24565
rect 42429 24565 42441 24599
rect 42475 24596 42487 24599
rect 43438 24596 43444 24608
rect 42475 24568 43444 24596
rect 42475 24565 42487 24568
rect 42429 24559 42487 24565
rect 43438 24556 43444 24568
rect 43496 24556 43502 24608
rect 44085 24599 44143 24605
rect 44085 24565 44097 24599
rect 44131 24596 44143 24599
rect 44910 24596 44916 24608
rect 44131 24568 44916 24596
rect 44131 24565 44143 24568
rect 44085 24559 44143 24565
rect 44910 24556 44916 24568
rect 44968 24556 44974 24608
rect 45388 24605 45416 24636
rect 45462 24624 45468 24676
rect 45520 24664 45526 24676
rect 46293 24667 46351 24673
rect 46293 24664 46305 24667
rect 45520 24636 46305 24664
rect 45520 24624 45526 24636
rect 46293 24633 46305 24636
rect 46339 24633 46351 24667
rect 46584 24664 46612 24772
rect 46661 24769 46673 24772
rect 46707 24769 46719 24803
rect 46661 24763 46719 24769
rect 46750 24760 46756 24812
rect 46808 24800 46814 24812
rect 46808 24772 46853 24800
rect 46808 24760 46814 24772
rect 47578 24760 47584 24812
rect 47636 24800 47642 24812
rect 47636 24772 47681 24800
rect 47636 24760 47642 24772
rect 56594 24760 56600 24812
rect 56652 24800 56658 24812
rect 56873 24803 56931 24809
rect 56873 24800 56885 24803
rect 56652 24772 56885 24800
rect 56652 24760 56658 24772
rect 56873 24769 56885 24772
rect 56919 24800 56931 24803
rect 57422 24800 57428 24812
rect 56919 24772 57428 24800
rect 56919 24769 56931 24772
rect 56873 24763 56931 24769
rect 57422 24760 57428 24772
rect 57480 24760 57486 24812
rect 47857 24735 47915 24741
rect 47857 24732 47869 24735
rect 47320 24704 47869 24732
rect 46658 24664 46664 24676
rect 46584 24636 46664 24664
rect 46293 24627 46351 24633
rect 46658 24624 46664 24636
rect 46716 24664 46722 24676
rect 47210 24664 47216 24676
rect 46716 24636 47216 24664
rect 46716 24624 46722 24636
rect 47210 24624 47216 24636
rect 47268 24624 47274 24676
rect 45373 24599 45431 24605
rect 45373 24565 45385 24599
rect 45419 24565 45431 24599
rect 45738 24596 45744 24608
rect 45699 24568 45744 24596
rect 45373 24559 45431 24565
rect 45738 24556 45744 24568
rect 45796 24556 45802 24608
rect 45830 24556 45836 24608
rect 45888 24596 45894 24608
rect 47320 24596 47348 24704
rect 47857 24701 47869 24704
rect 47903 24701 47915 24735
rect 47857 24695 47915 24701
rect 47946 24692 47952 24744
rect 48004 24732 48010 24744
rect 48004 24704 48049 24732
rect 48004 24692 48010 24704
rect 47578 24624 47584 24676
rect 47636 24664 47642 24676
rect 49234 24664 49240 24676
rect 47636 24636 49240 24664
rect 47636 24624 47642 24636
rect 49234 24624 49240 24636
rect 49292 24624 49298 24676
rect 47670 24596 47676 24608
rect 45888 24568 47348 24596
rect 47631 24568 47676 24596
rect 45888 24556 45894 24568
rect 47670 24556 47676 24568
rect 47728 24556 47734 24608
rect 56502 24556 56508 24608
rect 56560 24596 56566 24608
rect 56965 24599 57023 24605
rect 56965 24596 56977 24599
rect 56560 24568 56977 24596
rect 56560 24556 56566 24568
rect 56965 24565 56977 24568
rect 57011 24565 57023 24599
rect 58066 24596 58072 24608
rect 58027 24568 58072 24596
rect 56965 24559 57023 24565
rect 58066 24556 58072 24568
rect 58124 24556 58130 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 40310 24392 40316 24404
rect 40271 24364 40316 24392
rect 40310 24352 40316 24364
rect 40368 24352 40374 24404
rect 44453 24395 44511 24401
rect 44453 24361 44465 24395
rect 44499 24392 44511 24395
rect 44542 24392 44548 24404
rect 44499 24364 44548 24392
rect 44499 24361 44511 24364
rect 44453 24355 44511 24361
rect 44542 24352 44548 24364
rect 44600 24352 44606 24404
rect 46474 24352 46480 24404
rect 46532 24392 46538 24404
rect 46661 24395 46719 24401
rect 46661 24392 46673 24395
rect 46532 24364 46673 24392
rect 46532 24352 46538 24364
rect 46661 24361 46673 24364
rect 46707 24361 46719 24395
rect 46661 24355 46719 24361
rect 41966 24284 41972 24336
rect 42024 24324 42030 24336
rect 42794 24324 42800 24336
rect 42024 24296 42800 24324
rect 42024 24284 42030 24296
rect 42794 24284 42800 24296
rect 42852 24324 42858 24336
rect 43070 24324 43076 24336
rect 42852 24296 43076 24324
rect 42852 24284 42858 24296
rect 43070 24284 43076 24296
rect 43128 24324 43134 24336
rect 45830 24324 45836 24336
rect 43128 24296 45836 24324
rect 43128 24284 43134 24296
rect 45830 24284 45836 24296
rect 45888 24284 45894 24336
rect 46201 24327 46259 24333
rect 46201 24293 46213 24327
rect 46247 24324 46259 24327
rect 46934 24324 46940 24336
rect 46247 24296 46940 24324
rect 46247 24293 46259 24296
rect 46201 24287 46259 24293
rect 46934 24284 46940 24296
rect 46992 24324 46998 24336
rect 58066 24324 58072 24336
rect 46992 24296 48912 24324
rect 46992 24284 46998 24296
rect 32030 24216 32036 24268
rect 32088 24256 32094 24268
rect 32309 24259 32367 24265
rect 32309 24256 32321 24259
rect 32088 24228 32321 24256
rect 32088 24216 32094 24228
rect 32309 24225 32321 24228
rect 32355 24225 32367 24259
rect 40218 24256 40224 24268
rect 32309 24219 32367 24225
rect 39960 24228 40224 24256
rect 39298 24148 39304 24200
rect 39356 24188 39362 24200
rect 39960 24197 39988 24228
rect 40218 24216 40224 24228
rect 40276 24216 40282 24268
rect 41417 24259 41475 24265
rect 41417 24225 41429 24259
rect 41463 24256 41475 24259
rect 43993 24259 44051 24265
rect 41463 24228 43944 24256
rect 41463 24225 41475 24228
rect 41417 24219 41475 24225
rect 39945 24191 40003 24197
rect 39945 24188 39957 24191
rect 39356 24160 39957 24188
rect 39356 24148 39362 24160
rect 39945 24157 39957 24160
rect 39991 24157 40003 24191
rect 40126 24188 40132 24200
rect 40087 24160 40132 24188
rect 39945 24151 40003 24157
rect 40126 24148 40132 24160
rect 40184 24148 40190 24200
rect 41601 24191 41659 24197
rect 41601 24157 41613 24191
rect 41647 24188 41659 24191
rect 41690 24188 41696 24200
rect 41647 24160 41696 24188
rect 41647 24157 41659 24160
rect 41601 24151 41659 24157
rect 41690 24148 41696 24160
rect 41748 24148 41754 24200
rect 41874 24188 41880 24200
rect 41835 24160 41880 24188
rect 41874 24148 41880 24160
rect 41932 24148 41938 24200
rect 42705 24191 42763 24197
rect 42705 24157 42717 24191
rect 42751 24157 42763 24191
rect 42705 24151 42763 24157
rect 32493 24123 32551 24129
rect 32493 24089 32505 24123
rect 32539 24120 32551 24123
rect 32582 24120 32588 24132
rect 32539 24092 32588 24120
rect 32539 24089 32551 24092
rect 32493 24083 32551 24089
rect 32582 24080 32588 24092
rect 32640 24080 32646 24132
rect 34146 24120 34152 24132
rect 34107 24092 34152 24120
rect 34146 24080 34152 24092
rect 34204 24080 34210 24132
rect 41230 24080 41236 24132
rect 41288 24120 41294 24132
rect 41785 24123 41843 24129
rect 41785 24120 41797 24123
rect 41288 24092 41797 24120
rect 41288 24080 41294 24092
rect 41785 24089 41797 24092
rect 41831 24089 41843 24123
rect 41785 24083 41843 24089
rect 42720 24120 42748 24151
rect 42794 24148 42800 24200
rect 42852 24188 42858 24200
rect 42978 24188 42984 24200
rect 42852 24160 42897 24188
rect 42939 24160 42984 24188
rect 42852 24148 42858 24160
rect 42978 24148 42984 24160
rect 43036 24148 43042 24200
rect 42886 24120 42892 24132
rect 42720 24092 42892 24120
rect 41046 24012 41052 24064
rect 41104 24052 41110 24064
rect 42720 24052 42748 24092
rect 42886 24080 42892 24092
rect 42944 24120 42950 24132
rect 43622 24120 43628 24132
rect 42944 24092 43628 24120
rect 42944 24080 42950 24092
rect 43622 24080 43628 24092
rect 43680 24080 43686 24132
rect 43916 24120 43944 24228
rect 43993 24225 44005 24259
rect 44039 24256 44051 24259
rect 45738 24256 45744 24268
rect 44039 24228 45744 24256
rect 44039 24225 44051 24228
rect 43993 24219 44051 24225
rect 45738 24216 45744 24228
rect 45796 24216 45802 24268
rect 46290 24216 46296 24268
rect 46348 24256 46354 24268
rect 47213 24259 47271 24265
rect 47213 24256 47225 24259
rect 46348 24228 47225 24256
rect 46348 24216 46354 24228
rect 47213 24225 47225 24228
rect 47259 24225 47271 24259
rect 47946 24256 47952 24268
rect 47907 24228 47952 24256
rect 47213 24219 47271 24225
rect 47946 24216 47952 24228
rect 48004 24216 48010 24268
rect 44085 24191 44143 24197
rect 44085 24157 44097 24191
rect 44131 24188 44143 24191
rect 45186 24188 45192 24200
rect 44131 24160 45192 24188
rect 44131 24157 44143 24160
rect 44085 24151 44143 24157
rect 45186 24148 45192 24160
rect 45244 24148 45250 24200
rect 45922 24188 45928 24200
rect 45883 24160 45928 24188
rect 45922 24148 45928 24160
rect 45980 24148 45986 24200
rect 46017 24191 46075 24197
rect 46017 24157 46029 24191
rect 46063 24157 46075 24191
rect 46017 24151 46075 24157
rect 46032 24120 46060 24151
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 48884 24197 48912 24296
rect 56336 24296 58072 24324
rect 56336 24265 56364 24296
rect 58066 24284 58072 24296
rect 58124 24284 58130 24336
rect 56321 24259 56379 24265
rect 56321 24225 56333 24259
rect 56367 24225 56379 24259
rect 56502 24256 56508 24268
rect 56463 24228 56508 24256
rect 56321 24219 56379 24225
rect 56502 24216 56508 24228
rect 56560 24216 56566 24268
rect 58158 24256 58164 24268
rect 58119 24228 58164 24256
rect 58158 24216 58164 24228
rect 58216 24216 58222 24268
rect 48041 24191 48099 24197
rect 48041 24188 48053 24191
rect 47360 24160 48053 24188
rect 47360 24148 47366 24160
rect 48041 24157 48053 24160
rect 48087 24157 48099 24191
rect 48041 24151 48099 24157
rect 48869 24191 48927 24197
rect 48869 24157 48881 24191
rect 48915 24157 48927 24191
rect 48869 24151 48927 24157
rect 46566 24120 46572 24132
rect 43916 24092 46572 24120
rect 46566 24080 46572 24092
rect 46624 24080 46630 24132
rect 47029 24123 47087 24129
rect 47029 24089 47041 24123
rect 47075 24120 47087 24123
rect 49145 24123 49203 24129
rect 49145 24120 49157 24123
rect 47075 24092 49157 24120
rect 47075 24089 47087 24092
rect 47029 24083 47087 24089
rect 49145 24089 49157 24092
rect 49191 24089 49203 24123
rect 49145 24083 49203 24089
rect 41104 24024 42748 24052
rect 41104 24012 41110 24024
rect 44358 24012 44364 24064
rect 44416 24052 44422 24064
rect 45462 24052 45468 24064
rect 44416 24024 45468 24052
rect 44416 24012 44422 24024
rect 45462 24012 45468 24024
rect 45520 24012 45526 24064
rect 47121 24055 47179 24061
rect 47121 24021 47133 24055
rect 47167 24052 47179 24055
rect 48409 24055 48467 24061
rect 48409 24052 48421 24055
rect 47167 24024 48421 24052
rect 47167 24021 47179 24024
rect 47121 24015 47179 24021
rect 48409 24021 48421 24024
rect 48455 24021 48467 24055
rect 48409 24015 48467 24021
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 32582 23848 32588 23860
rect 32543 23820 32588 23848
rect 32582 23808 32588 23820
rect 32640 23808 32646 23860
rect 43625 23851 43683 23857
rect 43625 23817 43637 23851
rect 43671 23817 43683 23851
rect 43625 23811 43683 23817
rect 44085 23851 44143 23857
rect 44085 23817 44097 23851
rect 44131 23848 44143 23851
rect 44266 23848 44272 23860
rect 44131 23820 44272 23848
rect 44131 23817 44143 23820
rect 44085 23811 44143 23817
rect 2130 23780 2136 23792
rect 2091 23752 2136 23780
rect 2130 23740 2136 23752
rect 2188 23740 2194 23792
rect 43254 23740 43260 23792
rect 43312 23780 43318 23792
rect 43533 23783 43591 23789
rect 43533 23780 43545 23783
rect 43312 23752 43545 23780
rect 43312 23740 43318 23752
rect 43533 23749 43545 23752
rect 43579 23749 43591 23783
rect 43640 23780 43668 23811
rect 44266 23808 44272 23820
rect 44324 23808 44330 23860
rect 45186 23848 45192 23860
rect 45147 23820 45192 23848
rect 45186 23808 45192 23820
rect 45244 23808 45250 23860
rect 45462 23808 45468 23860
rect 45520 23848 45526 23860
rect 47946 23848 47952 23860
rect 45520 23820 47624 23848
rect 47907 23820 47952 23848
rect 45520 23808 45526 23820
rect 44453 23783 44511 23789
rect 44453 23780 44465 23783
rect 43640 23752 44465 23780
rect 43533 23743 43591 23749
rect 44453 23749 44465 23752
rect 44499 23780 44511 23783
rect 44499 23752 45600 23780
rect 44499 23749 44511 23752
rect 44453 23743 44511 23749
rect 1946 23712 1952 23724
rect 1907 23684 1952 23712
rect 1946 23672 1952 23684
rect 2004 23672 2010 23724
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23712 32551 23715
rect 33134 23712 33140 23724
rect 32539 23684 33140 23712
rect 32539 23681 32551 23684
rect 32493 23675 32551 23681
rect 33134 23672 33140 23684
rect 33192 23672 33198 23724
rect 43346 23712 43352 23724
rect 43307 23684 43352 23712
rect 43346 23672 43352 23684
rect 43404 23672 43410 23724
rect 43625 23715 43683 23721
rect 43625 23681 43637 23715
rect 43671 23712 43683 23715
rect 43806 23712 43812 23724
rect 43671 23684 43812 23712
rect 43671 23681 43683 23684
rect 43625 23675 43683 23681
rect 43806 23672 43812 23684
rect 43864 23672 43870 23724
rect 44269 23715 44327 23721
rect 44269 23681 44281 23715
rect 44315 23681 44327 23715
rect 44269 23675 44327 23681
rect 2774 23644 2780 23656
rect 2735 23616 2780 23644
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 44284 23588 44312 23675
rect 44358 23672 44364 23724
rect 44416 23712 44422 23724
rect 44634 23712 44640 23724
rect 44416 23684 44461 23712
rect 44595 23684 44640 23712
rect 44416 23672 44422 23684
rect 44634 23672 44640 23684
rect 44692 23672 44698 23724
rect 44726 23672 44732 23724
rect 44784 23712 44790 23724
rect 45462 23712 45468 23724
rect 44784 23684 44829 23712
rect 45423 23684 45468 23712
rect 44784 23672 44790 23684
rect 45462 23672 45468 23684
rect 45520 23672 45526 23724
rect 45572 23721 45600 23752
rect 46382 23740 46388 23792
rect 46440 23780 46446 23792
rect 47118 23780 47124 23792
rect 46440 23752 47124 23780
rect 46440 23740 46446 23752
rect 45557 23715 45615 23721
rect 45557 23681 45569 23715
rect 45603 23681 45615 23715
rect 45557 23675 45615 23681
rect 45922 23672 45928 23724
rect 45980 23712 45986 23724
rect 46658 23712 46664 23724
rect 45980 23684 46664 23712
rect 45980 23672 45986 23684
rect 46658 23672 46664 23684
rect 46716 23672 46722 23724
rect 46768 23721 46796 23752
rect 47118 23740 47124 23752
rect 47176 23740 47182 23792
rect 46753 23715 46811 23721
rect 46753 23681 46765 23715
rect 46799 23681 46811 23715
rect 46753 23675 46811 23681
rect 46845 23715 46903 23721
rect 46845 23681 46857 23715
rect 46891 23712 46903 23715
rect 47302 23712 47308 23724
rect 46891 23684 47308 23712
rect 46891 23681 46903 23684
rect 46845 23675 46903 23681
rect 47302 23672 47308 23684
rect 47360 23672 47366 23724
rect 47596 23721 47624 23820
rect 47946 23808 47952 23820
rect 48004 23808 48010 23860
rect 47581 23715 47639 23721
rect 47581 23681 47593 23715
rect 47627 23681 47639 23715
rect 47762 23712 47768 23724
rect 47723 23684 47768 23712
rect 47581 23675 47639 23681
rect 47762 23672 47768 23684
rect 47820 23672 47826 23724
rect 45373 23647 45431 23653
rect 45373 23613 45385 23647
rect 45419 23613 45431 23647
rect 45373 23607 45431 23613
rect 44266 23536 44272 23588
rect 44324 23576 44330 23588
rect 45388 23576 45416 23607
rect 45646 23604 45652 23656
rect 45704 23644 45710 23656
rect 46566 23644 46572 23656
rect 45704 23616 45749 23644
rect 46527 23616 46572 23644
rect 45704 23604 45710 23616
rect 46566 23604 46572 23616
rect 46624 23604 46630 23656
rect 46385 23579 46443 23585
rect 46385 23576 46397 23579
rect 44324 23548 46397 23576
rect 44324 23536 44330 23548
rect 46385 23545 46397 23548
rect 46431 23545 46443 23579
rect 46385 23539 46443 23545
rect 44634 23468 44640 23520
rect 44692 23508 44698 23520
rect 45646 23508 45652 23520
rect 44692 23480 45652 23508
rect 44692 23468 44698 23480
rect 45646 23468 45652 23480
rect 45704 23468 45710 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 43898 23264 43904 23316
rect 43956 23304 43962 23316
rect 45005 23307 45063 23313
rect 45005 23304 45017 23307
rect 43956 23276 45017 23304
rect 43956 23264 43962 23276
rect 45005 23273 45017 23276
rect 45051 23273 45063 23307
rect 45005 23267 45063 23273
rect 47029 23307 47087 23313
rect 47029 23273 47041 23307
rect 47075 23304 47087 23307
rect 47762 23304 47768 23316
rect 47075 23276 47768 23304
rect 47075 23273 47087 23276
rect 47029 23267 47087 23273
rect 47762 23264 47768 23276
rect 47820 23264 47826 23316
rect 40034 23196 40040 23248
rect 40092 23196 40098 23248
rect 40405 23239 40463 23245
rect 40405 23205 40417 23239
rect 40451 23236 40463 23239
rect 40451 23208 41000 23236
rect 40451 23205 40463 23208
rect 40405 23199 40463 23205
rect 40052 23168 40080 23196
rect 40972 23177 41000 23208
rect 40129 23171 40187 23177
rect 40129 23168 40141 23171
rect 40052 23140 40141 23168
rect 40129 23137 40141 23140
rect 40175 23137 40187 23171
rect 40129 23131 40187 23137
rect 40957 23171 41015 23177
rect 40957 23137 40969 23171
rect 41003 23137 41015 23171
rect 40957 23131 41015 23137
rect 41877 23171 41935 23177
rect 41877 23137 41889 23171
rect 41923 23168 41935 23171
rect 43254 23168 43260 23180
rect 41923 23140 43260 23168
rect 41923 23137 41935 23140
rect 41877 23131 41935 23137
rect 40037 23103 40095 23109
rect 40037 23069 40049 23103
rect 40083 23069 40095 23103
rect 40037 23063 40095 23069
rect 40052 22964 40080 23063
rect 40144 23032 40172 23131
rect 43254 23128 43260 23140
rect 43312 23128 43318 23180
rect 44085 23171 44143 23177
rect 44085 23137 44097 23171
rect 44131 23168 44143 23171
rect 44358 23168 44364 23180
rect 44131 23140 44364 23168
rect 44131 23137 44143 23140
rect 44085 23131 44143 23137
rect 44358 23128 44364 23140
rect 44416 23128 44422 23180
rect 45649 23171 45707 23177
rect 45649 23137 45661 23171
rect 45695 23168 45707 23171
rect 46290 23168 46296 23180
rect 45695 23140 46296 23168
rect 45695 23137 45707 23140
rect 45649 23131 45707 23137
rect 46290 23128 46296 23140
rect 46348 23128 46354 23180
rect 40402 23060 40408 23112
rect 40460 23100 40466 23112
rect 41049 23103 41107 23109
rect 41049 23100 41061 23103
rect 40460 23072 41061 23100
rect 40460 23060 40466 23072
rect 41049 23069 41061 23072
rect 41095 23069 41107 23103
rect 42061 23103 42119 23109
rect 42061 23100 42073 23103
rect 41049 23063 41107 23069
rect 41156 23072 42073 23100
rect 41156 23032 41184 23072
rect 42061 23069 42073 23072
rect 42107 23069 42119 23103
rect 42061 23063 42119 23069
rect 42337 23103 42395 23109
rect 42337 23069 42349 23103
rect 42383 23100 42395 23103
rect 42886 23100 42892 23112
rect 42383 23072 42892 23100
rect 42383 23069 42395 23072
rect 42337 23063 42395 23069
rect 42886 23060 42892 23072
rect 42944 23100 42950 23112
rect 42981 23103 43039 23109
rect 42981 23100 42993 23103
rect 42944 23072 42993 23100
rect 42944 23060 42950 23072
rect 42981 23069 42993 23072
rect 43027 23069 43039 23103
rect 42981 23063 43039 23069
rect 43070 23060 43076 23112
rect 43128 23100 43134 23112
rect 44266 23100 44272 23112
rect 43128 23072 43173 23100
rect 44227 23072 44272 23100
rect 43128 23060 43134 23072
rect 44266 23060 44272 23072
rect 44324 23060 44330 23112
rect 46934 23100 46940 23112
rect 46895 23072 46940 23100
rect 46934 23060 46940 23072
rect 46992 23060 46998 23112
rect 47118 23100 47124 23112
rect 47079 23072 47124 23100
rect 47118 23060 47124 23072
rect 47176 23060 47182 23112
rect 42797 23035 42855 23041
rect 42797 23032 42809 23035
rect 40144 23004 41184 23032
rect 41432 23004 42809 23032
rect 40678 22964 40684 22976
rect 40052 22936 40684 22964
rect 40678 22924 40684 22936
rect 40736 22924 40742 22976
rect 41432 22973 41460 23004
rect 42797 23001 42809 23004
rect 42843 23001 42855 23035
rect 43088 23032 43116 23060
rect 42797 22995 42855 23001
rect 42996 23004 43116 23032
rect 41417 22967 41475 22973
rect 41417 22933 41429 22967
rect 41463 22933 41475 22967
rect 41417 22927 41475 22933
rect 42245 22967 42303 22973
rect 42245 22933 42257 22967
rect 42291 22964 42303 22967
rect 42996 22964 43024 23004
rect 43714 22992 43720 23044
rect 43772 23032 43778 23044
rect 45373 23035 45431 23041
rect 45373 23032 45385 23035
rect 43772 23004 45385 23032
rect 43772 22992 43778 23004
rect 45373 23001 45385 23004
rect 45419 23001 45431 23035
rect 45373 22995 45431 23001
rect 42291 22936 43024 22964
rect 43073 22967 43131 22973
rect 42291 22933 42303 22936
rect 42245 22927 42303 22933
rect 43073 22933 43085 22967
rect 43119 22964 43131 22967
rect 43346 22964 43352 22976
rect 43119 22936 43352 22964
rect 43119 22933 43131 22936
rect 43073 22927 43131 22933
rect 43346 22924 43352 22936
rect 43404 22964 43410 22976
rect 43530 22964 43536 22976
rect 43404 22936 43536 22964
rect 43404 22924 43410 22936
rect 43530 22924 43536 22936
rect 43588 22924 43594 22976
rect 44358 22924 44364 22976
rect 44416 22964 44422 22976
rect 44453 22967 44511 22973
rect 44453 22964 44465 22967
rect 44416 22936 44465 22964
rect 44416 22924 44422 22936
rect 44453 22933 44465 22936
rect 44499 22933 44511 22967
rect 44453 22927 44511 22933
rect 45462 22924 45468 22976
rect 45520 22964 45526 22976
rect 45520 22936 45565 22964
rect 45520 22924 45526 22936
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 43714 22760 43720 22772
rect 43675 22732 43720 22760
rect 43714 22720 43720 22732
rect 43772 22720 43778 22772
rect 44729 22763 44787 22769
rect 44729 22729 44741 22763
rect 44775 22760 44787 22763
rect 45462 22760 45468 22772
rect 44775 22732 45468 22760
rect 44775 22729 44787 22732
rect 44729 22723 44787 22729
rect 45462 22720 45468 22732
rect 45520 22720 45526 22772
rect 57514 22692 57520 22704
rect 56520 22664 57520 22692
rect 43254 22584 43260 22636
rect 43312 22624 43318 22636
rect 43349 22627 43407 22633
rect 43349 22624 43361 22627
rect 43312 22596 43361 22624
rect 43312 22584 43318 22596
rect 43349 22593 43361 22596
rect 43395 22593 43407 22627
rect 43530 22624 43536 22636
rect 43491 22596 43536 22624
rect 43349 22587 43407 22593
rect 43530 22584 43536 22596
rect 43588 22584 43594 22636
rect 44358 22624 44364 22636
rect 44319 22596 44364 22624
rect 44358 22584 44364 22596
rect 44416 22584 44422 22636
rect 45186 22624 45192 22636
rect 45147 22596 45192 22624
rect 45186 22584 45192 22596
rect 45244 22584 45250 22636
rect 56520 22633 56548 22664
rect 57514 22652 57520 22664
rect 57572 22652 57578 22704
rect 45373 22627 45431 22633
rect 45373 22593 45385 22627
rect 45419 22593 45431 22627
rect 45373 22587 45431 22593
rect 56505 22627 56563 22633
rect 56505 22593 56517 22627
rect 56551 22593 56563 22627
rect 56505 22587 56563 22593
rect 57149 22627 57207 22633
rect 57149 22593 57161 22627
rect 57195 22624 57207 22627
rect 57606 22624 57612 22636
rect 57195 22596 57612 22624
rect 57195 22593 57207 22596
rect 57149 22587 57207 22593
rect 44453 22559 44511 22565
rect 44453 22525 44465 22559
rect 44499 22556 44511 22559
rect 45281 22559 45339 22565
rect 45281 22556 45293 22559
rect 44499 22528 45293 22556
rect 44499 22525 44511 22528
rect 44453 22519 44511 22525
rect 45281 22525 45293 22528
rect 45327 22525 45339 22559
rect 45281 22519 45339 22525
rect 44266 22448 44272 22500
rect 44324 22488 44330 22500
rect 45388 22488 45416 22587
rect 57606 22584 57612 22596
rect 57664 22584 57670 22636
rect 44324 22460 45416 22488
rect 44324 22448 44330 22460
rect 56594 22420 56600 22432
rect 56555 22392 56600 22420
rect 56594 22380 56600 22392
rect 56652 22380 56658 22432
rect 57238 22420 57244 22432
rect 57199 22392 57244 22420
rect 57238 22380 57244 22392
rect 57296 22380 57302 22432
rect 57330 22380 57336 22432
rect 57388 22420 57394 22432
rect 58069 22423 58127 22429
rect 58069 22420 58081 22423
rect 57388 22392 58081 22420
rect 57388 22380 57394 22392
rect 58069 22389 58081 22392
rect 58115 22389 58127 22423
rect 58069 22383 58127 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 43254 22176 43260 22228
rect 43312 22216 43318 22228
rect 43533 22219 43591 22225
rect 43533 22216 43545 22219
rect 43312 22188 43545 22216
rect 43312 22176 43318 22188
rect 43533 22185 43545 22188
rect 43579 22185 43591 22219
rect 43533 22179 43591 22185
rect 44177 22219 44235 22225
rect 44177 22185 44189 22219
rect 44223 22216 44235 22219
rect 44634 22216 44640 22228
rect 44223 22188 44640 22216
rect 44223 22185 44235 22188
rect 44177 22179 44235 22185
rect 43548 22148 43576 22179
rect 44634 22176 44640 22188
rect 44692 22216 44698 22228
rect 45186 22216 45192 22228
rect 44692 22188 45192 22216
rect 44692 22176 44698 22188
rect 45186 22176 45192 22188
rect 45244 22176 45250 22228
rect 57330 22148 57336 22160
rect 43548 22120 44128 22148
rect 43806 22080 43812 22092
rect 43364 22052 43812 22080
rect 1946 21972 1952 22024
rect 2004 22012 2010 22024
rect 2225 22015 2283 22021
rect 2225 22012 2237 22015
rect 2004 21984 2237 22012
rect 2004 21972 2010 21984
rect 2225 21981 2237 21984
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 43364 21953 43392 22052
rect 43806 22040 43812 22052
rect 43864 22040 43870 22092
rect 44100 22080 44128 22120
rect 56428 22120 57336 22148
rect 56321 22083 56379 22089
rect 44100 22052 44588 22080
rect 44453 22015 44511 22021
rect 44453 22012 44465 22015
rect 43640 21984 44465 22012
rect 43349 21947 43407 21953
rect 43349 21913 43361 21947
rect 43395 21913 43407 21947
rect 43530 21944 43536 21956
rect 43588 21953 43594 21956
rect 43588 21947 43612 21953
rect 43464 21916 43536 21944
rect 43349 21907 43407 21913
rect 43530 21904 43536 21916
rect 43600 21944 43612 21947
rect 43640 21944 43668 21984
rect 44453 21981 44465 21984
rect 44499 21981 44511 22015
rect 44453 21975 44511 21981
rect 43600 21916 43668 21944
rect 43600 21913 43612 21916
rect 43588 21907 43612 21913
rect 43588 21904 43594 21907
rect 43806 21904 43812 21956
rect 43864 21944 43870 21956
rect 44177 21947 44235 21953
rect 44177 21944 44189 21947
rect 43864 21916 44189 21944
rect 43864 21904 43870 21916
rect 44177 21913 44189 21916
rect 44223 21913 44235 21947
rect 44177 21907 44235 21913
rect 43717 21879 43775 21885
rect 43717 21845 43729 21879
rect 43763 21876 43775 21879
rect 44266 21876 44272 21888
rect 43763 21848 44272 21876
rect 43763 21845 43775 21848
rect 43717 21839 43775 21845
rect 44266 21836 44272 21848
rect 44324 21836 44330 21888
rect 44361 21879 44419 21885
rect 44361 21845 44373 21879
rect 44407 21876 44419 21879
rect 44560 21876 44588 22052
rect 56321 22049 56333 22083
rect 56367 22080 56379 22083
rect 56428 22080 56456 22120
rect 57330 22108 57336 22120
rect 57388 22108 57394 22160
rect 56367 22052 56456 22080
rect 56505 22083 56563 22089
rect 56367 22049 56379 22052
rect 56321 22043 56379 22049
rect 56505 22049 56517 22083
rect 56551 22080 56563 22083
rect 56594 22080 56600 22092
rect 56551 22052 56600 22080
rect 56551 22049 56563 22052
rect 56505 22043 56563 22049
rect 56594 22040 56600 22052
rect 56652 22040 56658 22092
rect 57882 22080 57888 22092
rect 57843 22052 57888 22080
rect 57882 22040 57888 22052
rect 57940 22040 57946 22092
rect 44407 21848 44588 21876
rect 44407 21845 44419 21848
rect 44361 21839 44419 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 17126 21672 17132 21684
rect 17087 21644 17132 21672
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 1946 21536 1952 21548
rect 1907 21508 1952 21536
rect 1946 21496 1952 21508
rect 2004 21496 2010 21548
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21536 17095 21539
rect 17402 21536 17408 21548
rect 17083 21508 17408 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 17402 21496 17408 21508
rect 17460 21496 17466 21548
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19613 21539 19671 21545
rect 19613 21536 19625 21539
rect 19484 21508 19625 21536
rect 19484 21496 19490 21508
rect 19613 21505 19625 21508
rect 19659 21505 19671 21539
rect 19613 21499 19671 21505
rect 29638 21496 29644 21548
rect 29696 21536 29702 21548
rect 29733 21539 29791 21545
rect 29733 21536 29745 21539
rect 29696 21508 29745 21536
rect 29696 21496 29702 21508
rect 29733 21505 29745 21508
rect 29779 21505 29791 21539
rect 56965 21539 57023 21545
rect 56965 21536 56977 21539
rect 29733 21499 29791 21505
rect 45526 21508 56977 21536
rect 2130 21468 2136 21480
rect 2091 21440 2136 21468
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 2774 21468 2780 21480
rect 2735 21440 2780 21468
rect 2774 21428 2780 21440
rect 2832 21428 2838 21480
rect 20165 21471 20223 21477
rect 20165 21437 20177 21471
rect 20211 21468 20223 21471
rect 20254 21468 20260 21480
rect 20211 21440 20260 21468
rect 20211 21437 20223 21440
rect 20165 21431 20223 21437
rect 20254 21428 20260 21440
rect 20312 21428 20318 21480
rect 31481 21471 31539 21477
rect 31481 21437 31493 21471
rect 31527 21437 31539 21471
rect 31481 21431 31539 21437
rect 31496 21400 31524 21431
rect 45526 21400 45554 21508
rect 56965 21505 56977 21508
rect 57011 21536 57023 21539
rect 57698 21536 57704 21548
rect 57011 21508 57704 21536
rect 57011 21505 57023 21508
rect 56965 21499 57023 21505
rect 57698 21496 57704 21508
rect 57756 21496 57762 21548
rect 26206 21372 45554 21400
rect 3878 21292 3884 21344
rect 3936 21332 3942 21344
rect 26206 21332 26234 21372
rect 57054 21332 57060 21344
rect 3936 21304 26234 21332
rect 57015 21304 57060 21332
rect 3936 21292 3942 21304
rect 57054 21292 57060 21304
rect 57112 21292 57118 21344
rect 57146 21292 57152 21344
rect 57204 21332 57210 21344
rect 58069 21335 58127 21341
rect 58069 21332 58081 21335
rect 57204 21304 58081 21332
rect 57204 21292 57210 21304
rect 58069 21301 58081 21304
rect 58115 21301 58127 21335
rect 58069 21295 58127 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 18432 20964 26234 20992
rect 1946 20884 1952 20936
rect 2004 20924 2010 20936
rect 18432 20933 18460 20964
rect 2225 20927 2283 20933
rect 2225 20924 2237 20927
rect 2004 20896 2237 20924
rect 2004 20884 2010 20896
rect 2225 20893 2237 20896
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20893 18475 20927
rect 19426 20924 19432 20936
rect 18417 20887 18475 20893
rect 18616 20896 19432 20924
rect 18616 20797 18644 20896
rect 19426 20884 19432 20896
rect 19484 20924 19490 20936
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19484 20896 19625 20924
rect 19484 20884 19490 20896
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 26206 20924 26234 20964
rect 31202 20952 31208 21004
rect 31260 20992 31266 21004
rect 31297 20995 31355 21001
rect 31297 20992 31309 20995
rect 31260 20964 31309 20992
rect 31260 20952 31266 20964
rect 31297 20961 31309 20964
rect 31343 20992 31355 20995
rect 35342 20992 35348 21004
rect 31343 20964 35348 20992
rect 31343 20961 31355 20964
rect 31297 20955 31355 20961
rect 35342 20952 35348 20964
rect 35400 20952 35406 21004
rect 56321 20995 56379 21001
rect 56321 20961 56333 20995
rect 56367 20992 56379 20995
rect 57882 20992 57888 21004
rect 56367 20964 57744 20992
rect 57843 20964 57888 20992
rect 56367 20961 56379 20964
rect 56321 20955 56379 20961
rect 28442 20924 28448 20936
rect 26206 20896 28448 20924
rect 19613 20887 19671 20893
rect 28442 20884 28448 20896
rect 28500 20924 28506 20936
rect 28629 20927 28687 20933
rect 28629 20924 28641 20927
rect 28500 20896 28641 20924
rect 28500 20884 28506 20896
rect 28629 20893 28641 20896
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 30469 20927 30527 20933
rect 30469 20893 30481 20927
rect 30515 20893 30527 20927
rect 57716 20924 57744 20964
rect 57882 20952 57888 20964
rect 57940 20952 57946 21004
rect 58066 20924 58072 20936
rect 57716 20896 58072 20924
rect 30469 20887 30527 20893
rect 20165 20859 20223 20865
rect 20165 20825 20177 20859
rect 20211 20825 20223 20859
rect 20165 20819 20223 20825
rect 28997 20859 29055 20865
rect 28997 20825 29009 20859
rect 29043 20856 29055 20859
rect 29638 20856 29644 20868
rect 29043 20828 29644 20856
rect 29043 20825 29055 20828
rect 28997 20819 29055 20825
rect 18601 20791 18659 20797
rect 18601 20757 18613 20791
rect 18647 20757 18659 20791
rect 18601 20751 18659 20757
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 20180 20788 20208 20819
rect 29638 20816 29644 20828
rect 29696 20856 29702 20868
rect 30484 20856 30512 20887
rect 58066 20884 58072 20896
rect 58124 20884 58130 20936
rect 29696 20828 30512 20856
rect 56505 20859 56563 20865
rect 29696 20816 29702 20828
rect 56505 20825 56517 20859
rect 56551 20856 56563 20859
rect 57238 20856 57244 20868
rect 56551 20828 57244 20856
rect 56551 20825 56563 20828
rect 56505 20819 56563 20825
rect 57238 20816 57244 20828
rect 57296 20816 57302 20868
rect 47578 20788 47584 20800
rect 19392 20760 47584 20788
rect 19392 20748 19398 20760
rect 47578 20748 47584 20760
rect 47636 20748 47642 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 30466 20476 30472 20528
rect 30524 20516 30530 20528
rect 30561 20519 30619 20525
rect 30561 20516 30573 20519
rect 30524 20488 30573 20516
rect 30524 20476 30530 20488
rect 30561 20485 30573 20488
rect 30607 20485 30619 20519
rect 30561 20479 30619 20485
rect 1946 20448 1952 20460
rect 1907 20420 1952 20448
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 19521 20451 19579 20457
rect 19521 20448 19533 20451
rect 19484 20420 19533 20448
rect 19484 20408 19490 20420
rect 19521 20417 19533 20420
rect 19567 20417 19579 20451
rect 29638 20448 29644 20460
rect 29599 20420 29644 20448
rect 19521 20411 19579 20417
rect 29638 20408 29644 20420
rect 29696 20408 29702 20460
rect 58066 20448 58072 20460
rect 58027 20420 58072 20448
rect 58066 20408 58072 20420
rect 58124 20408 58130 20460
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20380 2191 20383
rect 2498 20380 2504 20392
rect 2179 20352 2504 20380
rect 2179 20349 2191 20352
rect 2133 20343 2191 20349
rect 2498 20340 2504 20352
rect 2556 20340 2562 20392
rect 2774 20380 2780 20392
rect 2735 20352 2780 20380
rect 2774 20340 2780 20352
rect 2832 20340 2838 20392
rect 3970 20340 3976 20392
rect 4028 20380 4034 20392
rect 20346 20380 20352 20392
rect 4028 20352 20352 20380
rect 4028 20340 4034 20352
rect 20346 20340 20352 20352
rect 20404 20340 20410 20392
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 2130 20000 2136 20052
rect 2188 20040 2194 20052
rect 2593 20043 2651 20049
rect 2593 20040 2605 20043
rect 2188 20012 2605 20040
rect 2188 20000 2194 20012
rect 2593 20009 2605 20012
rect 2639 20009 2651 20043
rect 2593 20003 2651 20009
rect 57146 19972 57152 19984
rect 56336 19944 57152 19972
rect 31110 19904 31116 19916
rect 31071 19876 31116 19904
rect 31110 19864 31116 19876
rect 31168 19904 31174 19916
rect 56336 19913 56364 19944
rect 57146 19932 57152 19944
rect 57204 19932 57210 19984
rect 56321 19907 56379 19913
rect 31168 19876 35894 19904
rect 31168 19864 31174 19876
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19836 2559 19839
rect 2682 19836 2688 19848
rect 2547 19808 2688 19836
rect 2547 19805 2559 19808
rect 2501 19799 2559 19805
rect 2682 19796 2688 19808
rect 2740 19836 2746 19848
rect 19334 19836 19340 19848
rect 2740 19808 19340 19836
rect 2740 19796 2746 19808
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 19426 19796 19432 19848
rect 19484 19836 19490 19848
rect 19521 19839 19579 19845
rect 19521 19836 19533 19839
rect 19484 19808 19533 19836
rect 19484 19796 19490 19808
rect 19521 19805 19533 19808
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 29638 19796 29644 19848
rect 29696 19836 29702 19848
rect 30469 19839 30527 19845
rect 30469 19836 30481 19839
rect 29696 19808 30481 19836
rect 29696 19796 29702 19808
rect 30469 19805 30481 19808
rect 30515 19805 30527 19839
rect 30469 19799 30527 19805
rect 12434 19728 12440 19780
rect 12492 19768 12498 19780
rect 12986 19768 12992 19780
rect 12492 19740 12992 19768
rect 12492 19728 12498 19740
rect 12986 19728 12992 19740
rect 13044 19768 13050 19780
rect 20438 19768 20444 19780
rect 13044 19740 20444 19768
rect 13044 19728 13050 19740
rect 20438 19728 20444 19740
rect 20496 19728 20502 19780
rect 35866 19768 35894 19876
rect 56321 19873 56333 19907
rect 56367 19873 56379 19907
rect 56321 19867 56379 19873
rect 56505 19907 56563 19913
rect 56505 19873 56517 19907
rect 56551 19904 56563 19907
rect 57054 19904 57060 19916
rect 56551 19876 57060 19904
rect 56551 19873 56563 19876
rect 56505 19867 56563 19873
rect 57054 19864 57060 19876
rect 57112 19864 57118 19916
rect 57790 19904 57796 19916
rect 57751 19876 57796 19904
rect 57790 19864 57796 19876
rect 57848 19864 57854 19916
rect 46750 19768 46756 19780
rect 35866 19740 46756 19768
rect 46750 19728 46756 19740
rect 46808 19728 46814 19780
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 2498 19496 2504 19508
rect 2459 19468 2504 19496
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 2406 19360 2412 19372
rect 2367 19332 2412 19360
rect 2406 19320 2412 19332
rect 2464 19360 2470 19372
rect 12434 19360 12440 19372
rect 2464 19332 12440 19360
rect 2464 19320 2470 19332
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19484 19332 19533 19360
rect 19484 19320 19490 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 20070 19360 20076 19372
rect 20031 19332 20076 19360
rect 19521 19323 19579 19329
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 29549 19363 29607 19369
rect 29549 19329 29561 19363
rect 29595 19360 29607 19363
rect 29638 19360 29644 19372
rect 29595 19332 29644 19360
rect 29595 19329 29607 19332
rect 29549 19323 29607 19329
rect 29638 19320 29644 19332
rect 29696 19320 29702 19372
rect 29825 19363 29883 19369
rect 29825 19329 29837 19363
rect 29871 19360 29883 19363
rect 30374 19360 30380 19372
rect 29871 19332 30380 19360
rect 29871 19329 29883 19332
rect 29825 19323 29883 19329
rect 30374 19320 30380 19332
rect 30432 19320 30438 19372
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 2501 18751 2559 18757
rect 2501 18748 2513 18751
rect 2280 18720 2513 18748
rect 2280 18708 2286 18720
rect 2501 18717 2513 18720
rect 2547 18717 2559 18751
rect 2501 18711 2559 18717
rect 3789 18751 3847 18757
rect 3789 18717 3801 18751
rect 3835 18748 3847 18751
rect 9030 18748 9036 18760
rect 3835 18720 9036 18748
rect 3835 18717 3847 18720
rect 3789 18711 3847 18717
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 2406 18572 2412 18624
rect 2464 18612 2470 18624
rect 3881 18615 3939 18621
rect 3881 18612 3893 18615
rect 2464 18584 3893 18612
rect 2464 18572 2470 18584
rect 3881 18581 3893 18584
rect 3927 18581 3939 18615
rect 3881 18575 3939 18581
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 2406 18340 2412 18352
rect 2367 18312 2412 18340
rect 2406 18300 2412 18312
rect 2464 18300 2470 18352
rect 2222 18272 2228 18284
rect 2183 18244 2228 18272
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 30374 18272 30380 18284
rect 30335 18244 30380 18272
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 2774 18204 2780 18216
rect 2735 18176 2780 18204
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 30469 18071 30527 18077
rect 30469 18037 30481 18071
rect 30515 18068 30527 18071
rect 31202 18068 31208 18080
rect 30515 18040 31208 18068
rect 30515 18037 30527 18040
rect 30469 18031 30527 18037
rect 31202 18028 31208 18040
rect 31260 18028 31266 18080
rect 56870 18028 56876 18080
rect 56928 18068 56934 18080
rect 58069 18071 58127 18077
rect 58069 18068 58081 18071
rect 56928 18040 58081 18068
rect 56928 18028 56934 18040
rect 58069 18037 58081 18040
rect 58115 18037 58127 18071
rect 58069 18031 58127 18037
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 31018 17728 31024 17740
rect 30979 17700 31024 17728
rect 31018 17688 31024 17700
rect 31076 17688 31082 17740
rect 31202 17728 31208 17740
rect 31163 17700 31208 17728
rect 31202 17688 31208 17700
rect 31260 17688 31266 17740
rect 56321 17731 56379 17737
rect 56321 17697 56333 17731
rect 56367 17728 56379 17731
rect 56870 17728 56876 17740
rect 56367 17700 56876 17728
rect 56367 17697 56379 17700
rect 56321 17691 56379 17697
rect 56870 17688 56876 17700
rect 56928 17688 56934 17740
rect 58158 17728 58164 17740
rect 58119 17700 58164 17728
rect 58158 17688 58164 17700
rect 58216 17688 58222 17740
rect 1946 17620 1952 17672
rect 2004 17660 2010 17672
rect 2225 17663 2283 17669
rect 2225 17660 2237 17663
rect 2004 17632 2237 17660
rect 2004 17620 2010 17632
rect 2225 17629 2237 17632
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 32858 17592 32864 17604
rect 32819 17564 32864 17592
rect 32858 17552 32864 17564
rect 32916 17552 32922 17604
rect 56505 17595 56563 17601
rect 56505 17561 56517 17595
rect 56551 17592 56563 17595
rect 57146 17592 57152 17604
rect 56551 17564 57152 17592
rect 56551 17561 56563 17564
rect 56505 17555 56563 17561
rect 57146 17552 57152 17564
rect 57204 17552 57210 17604
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 57146 17320 57152 17332
rect 57107 17292 57152 17320
rect 57146 17280 57152 17292
rect 57204 17280 57210 17332
rect 1946 17184 1952 17196
rect 1907 17156 1952 17184
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 17402 17144 17408 17196
rect 17460 17184 17466 17196
rect 20070 17184 20076 17196
rect 17460 17156 20076 17184
rect 17460 17144 17466 17156
rect 20070 17144 20076 17156
rect 20128 17184 20134 17196
rect 57054 17184 57060 17196
rect 20128 17156 57060 17184
rect 20128 17144 20134 17156
rect 57054 17144 57060 17156
rect 57112 17144 57118 17196
rect 2130 17116 2136 17128
rect 2091 17088 2136 17116
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 56318 16940 56324 16992
rect 56376 16980 56382 16992
rect 58069 16983 58127 16989
rect 58069 16980 58081 16983
rect 56376 16952 58081 16980
rect 56376 16940 56382 16952
rect 58069 16949 58081 16952
rect 58115 16949 58127 16983
rect 58069 16943 58127 16949
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 2130 16736 2136 16788
rect 2188 16776 2194 16788
rect 2409 16779 2467 16785
rect 2409 16776 2421 16779
rect 2188 16748 2421 16776
rect 2188 16736 2194 16748
rect 2409 16745 2421 16748
rect 2455 16745 2467 16779
rect 2409 16739 2467 16745
rect 2038 16600 2044 16652
rect 2096 16640 2102 16652
rect 29546 16640 29552 16652
rect 2096 16612 29552 16640
rect 2096 16600 2102 16612
rect 2332 16581 2360 16612
rect 29546 16600 29552 16612
rect 29604 16640 29610 16652
rect 30282 16640 30288 16652
rect 29604 16612 30288 16640
rect 29604 16600 29610 16612
rect 30282 16600 30288 16612
rect 30340 16600 30346 16652
rect 56318 16640 56324 16652
rect 56279 16612 56324 16640
rect 56318 16600 56324 16612
rect 56376 16600 56382 16652
rect 57790 16640 57796 16652
rect 57751 16612 57796 16640
rect 57790 16600 57796 16612
rect 57848 16600 57854 16652
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16574 2375 16575
rect 2363 16546 2397 16574
rect 2363 16541 2375 16546
rect 2317 16535 2375 16541
rect 56505 16507 56563 16513
rect 56505 16473 56517 16507
rect 56551 16504 56563 16507
rect 57146 16504 57152 16516
rect 56551 16476 57152 16504
rect 56551 16473 56563 16476
rect 56505 16467 56563 16473
rect 57146 16464 57152 16476
rect 57204 16464 57210 16516
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 57146 16232 57152 16244
rect 57107 16204 57152 16232
rect 57146 16192 57152 16204
rect 57204 16192 57210 16244
rect 57054 16096 57060 16108
rect 57015 16068 57060 16096
rect 57054 16056 57060 16068
rect 57112 16056 57118 16108
rect 56318 15852 56324 15904
rect 56376 15892 56382 15904
rect 58069 15895 58127 15901
rect 58069 15892 58081 15895
rect 56376 15864 58081 15892
rect 56376 15852 56382 15864
rect 58069 15861 58081 15864
rect 58115 15861 58127 15895
rect 58069 15855 58127 15861
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 56318 15552 56324 15564
rect 56279 15524 56324 15552
rect 56318 15512 56324 15524
rect 56376 15512 56382 15564
rect 57882 15552 57888 15564
rect 57843 15524 57888 15552
rect 57882 15512 57888 15524
rect 57940 15512 57946 15564
rect 56505 15419 56563 15425
rect 56505 15385 56517 15419
rect 56551 15416 56563 15419
rect 56962 15416 56968 15428
rect 56551 15388 56968 15416
rect 56551 15385 56563 15388
rect 56505 15379 56563 15385
rect 56962 15376 56968 15388
rect 57020 15376 57026 15428
rect 57054 15308 57060 15360
rect 57112 15348 57118 15360
rect 57790 15348 57796 15360
rect 57112 15320 57796 15348
rect 57112 15308 57118 15320
rect 57790 15308 57796 15320
rect 57848 15308 57854 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 56962 15144 56968 15156
rect 56923 15116 56968 15144
rect 56962 15104 56968 15116
rect 57020 15104 57026 15156
rect 55674 14968 55680 15020
rect 55732 15008 55738 15020
rect 56873 15011 56931 15017
rect 56873 15008 56885 15011
rect 55732 14980 56885 15008
rect 55732 14968 55738 14980
rect 56873 14977 56885 14980
rect 56919 15008 56931 15011
rect 57330 15008 57336 15020
rect 56919 14980 57336 15008
rect 56919 14977 56931 14980
rect 56873 14971 56931 14977
rect 57330 14968 57336 14980
rect 57388 14968 57394 15020
rect 56318 14764 56324 14816
rect 56376 14804 56382 14816
rect 58069 14807 58127 14813
rect 58069 14804 58081 14807
rect 56376 14776 58081 14804
rect 56376 14764 56382 14776
rect 58069 14773 58081 14776
rect 58115 14773 58127 14807
rect 58069 14767 58127 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 56318 14464 56324 14476
rect 56279 14436 56324 14464
rect 56318 14424 56324 14436
rect 56376 14424 56382 14476
rect 1946 14356 1952 14408
rect 2004 14396 2010 14408
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 2004 14368 2237 14396
rect 2004 14356 2010 14368
rect 2225 14365 2237 14368
rect 2271 14365 2283 14399
rect 2225 14359 2283 14365
rect 56505 14331 56563 14337
rect 56505 14297 56517 14331
rect 56551 14328 56563 14331
rect 56962 14328 56968 14340
rect 56551 14300 56968 14328
rect 56551 14297 56563 14300
rect 56505 14291 56563 14297
rect 56962 14288 56968 14300
rect 57020 14288 57026 14340
rect 58158 14328 58164 14340
rect 58119 14300 58164 14328
rect 58158 14288 58164 14300
rect 58216 14288 58222 14340
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 56962 14056 56968 14068
rect 56923 14028 56968 14056
rect 56962 14016 56968 14028
rect 57020 14016 57026 14068
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 56873 13923 56931 13929
rect 56873 13889 56885 13923
rect 56919 13920 56931 13923
rect 57146 13920 57152 13932
rect 56919 13892 57152 13920
rect 56919 13889 56931 13892
rect 56873 13883 56931 13889
rect 57146 13880 57152 13892
rect 57204 13880 57210 13932
rect 2130 13852 2136 13864
rect 2091 13824 2136 13852
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2774 13852 2780 13864
rect 2735 13824 2780 13852
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 2130 13472 2136 13524
rect 2188 13512 2194 13524
rect 2501 13515 2559 13521
rect 2501 13512 2513 13515
rect 2188 13484 2513 13512
rect 2188 13472 2194 13484
rect 2501 13481 2513 13484
rect 2547 13481 2559 13515
rect 2501 13475 2559 13481
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2682 13308 2688 13320
rect 2455 13280 2688 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2682 13268 2688 13280
rect 2740 13308 2746 13320
rect 4706 13308 4712 13320
rect 2740 13280 4712 13308
rect 2740 13268 2746 13280
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 2225 12767 2283 12773
rect 2225 12764 2237 12767
rect 1811 12736 2237 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 2225 12733 2237 12736
rect 2271 12733 2283 12767
rect 2225 12727 2283 12733
rect 2409 12767 2467 12773
rect 2409 12733 2421 12767
rect 2455 12764 2467 12767
rect 3878 12764 3884 12776
rect 2455 12736 3884 12764
rect 2455 12733 2467 12736
rect 2409 12727 2467 12733
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 4028 12736 4073 12764
rect 4028 12724 4034 12736
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 3878 12424 3884 12436
rect 3839 12396 3884 12424
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 2004 12192 2237 12220
rect 2004 12180 2010 12192
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12220 3847 12223
rect 14826 12220 14832 12232
rect 3835 12192 14832 12220
rect 3835 12189 3847 12192
rect 3789 12183 3847 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2406 11676 2412 11688
rect 2179 11648 2412 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 2406 11336 2412 11348
rect 2367 11308 2412 11336
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11132 2378 11144
rect 9122 11132 9128 11144
rect 2372 11104 9128 11132
rect 2372 11092 2378 11104
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 20346 10140 20352 10192
rect 20404 10180 20410 10192
rect 56686 10180 56692 10192
rect 20404 10152 56692 10180
rect 20404 10140 20410 10152
rect 56686 10140 56692 10152
rect 56744 10140 56750 10192
rect 30009 10115 30067 10121
rect 30009 10112 30021 10115
rect 26206 10084 30021 10112
rect 3418 9936 3424 9988
rect 3476 9976 3482 9988
rect 26206 9976 26234 10084
rect 30009 10081 30021 10084
rect 30055 10081 30067 10115
rect 57977 10115 58035 10121
rect 57977 10112 57989 10115
rect 30009 10075 30067 10081
rect 35866 10084 57989 10112
rect 29362 10004 29368 10056
rect 29420 10044 29426 10056
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 29420 10016 29561 10044
rect 29420 10004 29426 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29549 10007 29607 10013
rect 29730 9976 29736 9988
rect 3476 9948 26234 9976
rect 29691 9948 29736 9976
rect 3476 9936 3482 9948
rect 29730 9936 29736 9948
rect 29788 9936 29794 9988
rect 27154 9868 27160 9920
rect 27212 9908 27218 9920
rect 35866 9908 35894 10084
rect 57977 10081 57989 10084
rect 58023 10081 58035 10115
rect 57977 10075 58035 10081
rect 56597 10047 56655 10053
rect 56597 10013 56609 10047
rect 56643 10044 56655 10047
rect 56686 10044 56692 10056
rect 56643 10016 56692 10044
rect 56643 10013 56655 10016
rect 56597 10007 56655 10013
rect 56686 10004 56692 10016
rect 56744 10004 56750 10056
rect 57238 9976 57244 9988
rect 57199 9948 57244 9976
rect 57238 9936 57244 9948
rect 57296 9936 57302 9988
rect 56686 9908 56692 9920
rect 27212 9880 35894 9908
rect 56647 9880 56692 9908
rect 27212 9868 27218 9880
rect 56686 9868 56692 9880
rect 56744 9868 56750 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 29641 9707 29699 9713
rect 29641 9673 29653 9707
rect 29687 9704 29699 9707
rect 29730 9704 29736 9716
rect 29687 9676 29736 9704
rect 29687 9673 29699 9676
rect 29641 9667 29699 9673
rect 29730 9664 29736 9676
rect 29788 9664 29794 9716
rect 29546 9568 29552 9580
rect 29507 9540 29552 9568
rect 29546 9528 29552 9540
rect 29604 9528 29610 9580
rect 56318 9324 56324 9376
rect 56376 9364 56382 9376
rect 58069 9367 58127 9373
rect 58069 9364 58081 9367
rect 56376 9336 58081 9364
rect 56376 9324 56382 9336
rect 58069 9333 58081 9336
rect 58115 9333 58127 9367
rect 58069 9327 58127 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 56318 9024 56324 9036
rect 56279 8996 56324 9024
rect 56318 8984 56324 8996
rect 56376 8984 56382 9036
rect 56505 9027 56563 9033
rect 56505 8993 56517 9027
rect 56551 9024 56563 9027
rect 56686 9024 56692 9036
rect 56551 8996 56692 9024
rect 56551 8993 56563 8996
rect 56505 8987 56563 8993
rect 56686 8984 56692 8996
rect 56744 8984 56750 9036
rect 57882 9024 57888 9036
rect 57843 8996 57888 9024
rect 57882 8984 57888 8996
rect 57940 8984 57946 9036
rect 1946 8916 1952 8968
rect 2004 8956 2010 8968
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 2004 8928 2237 8956
rect 2004 8916 2010 8928
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2130 8412 2136 8424
rect 2091 8384 2136 8412
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2774 8412 2780 8424
rect 2735 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 2130 8072 2136 8084
rect 2091 8044 2136 8072
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1946 7868 1952 7880
rect 1627 7840 1952 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2685 7871 2743 7877
rect 2096 7840 2141 7868
rect 2096 7828 2102 7840
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 9858 7868 9864 7880
rect 2731 7840 9864 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 2777 7735 2835 7741
rect 2777 7732 2789 7735
rect 2188 7704 2789 7732
rect 2188 7692 2194 7704
rect 2777 7701 2789 7704
rect 2823 7701 2835 7735
rect 2777 7695 2835 7701
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 2130 7460 2136 7472
rect 2091 7432 2136 7460
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 20254 7392 20260 7404
rect 4295 7364 20260 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 2774 7324 2780 7336
rect 2735 7296 2780 7324
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4614 7188 4620 7200
rect 4387 7160 4620 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 1443 6820 3985 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 4614 6780 4620 6792
rect 3160 6752 4620 6780
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 3160 6712 3188 6752
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 56870 6780 56876 6792
rect 20496 6752 56876 6780
rect 20496 6740 20502 6752
rect 56870 6740 56876 6752
rect 56928 6780 56934 6792
rect 56965 6783 57023 6789
rect 56965 6780 56977 6783
rect 56928 6752 56977 6780
rect 56928 6740 56934 6752
rect 56965 6749 56977 6752
rect 57011 6749 57023 6783
rect 56965 6743 57023 6749
rect 57793 6783 57851 6789
rect 57793 6749 57805 6783
rect 57839 6749 57851 6783
rect 57793 6743 57851 6749
rect 1627 6684 3188 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 3292 6684 3337 6712
rect 3292 6672 3298 6684
rect 56318 6672 56324 6724
rect 56376 6712 56382 6724
rect 57808 6712 57836 6743
rect 56376 6684 57836 6712
rect 56376 6672 56382 6684
rect 57054 6644 57060 6656
rect 57015 6616 57060 6644
rect 57054 6604 57060 6616
rect 57112 6604 57118 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 5166 6372 5172 6384
rect 3016 6344 4292 6372
rect 5127 6344 5172 6372
rect 3016 6332 3022 6344
rect 4264 6313 4292 6344
rect 5166 6332 5172 6344
rect 5224 6372 5230 6384
rect 7834 6372 7840 6384
rect 5224 6344 7840 6372
rect 5224 6332 5230 6344
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 29454 6264 29460 6316
rect 29512 6304 29518 6316
rect 55585 6307 55643 6313
rect 55585 6304 55597 6307
rect 29512 6276 55597 6304
rect 29512 6264 29518 6276
rect 55585 6273 55597 6276
rect 55631 6304 55643 6307
rect 57885 6307 57943 6313
rect 57885 6304 57897 6307
rect 55631 6276 57897 6304
rect 55631 6273 55643 6276
rect 55585 6267 55643 6273
rect 57885 6273 57897 6276
rect 57931 6273 57943 6307
rect 57885 6267 57943 6273
rect 1854 6196 1860 6248
rect 1912 6236 1918 6248
rect 1949 6239 2007 6245
rect 1949 6236 1961 6239
rect 1912 6208 1961 6236
rect 1912 6196 1918 6208
rect 1949 6205 1961 6208
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6236 2191 6239
rect 2406 6236 2412 6248
rect 2179 6208 2412 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2866 6236 2872 6248
rect 2827 6208 2872 6236
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 56594 6060 56600 6112
rect 56652 6100 56658 6112
rect 56873 6103 56931 6109
rect 56873 6100 56885 6103
rect 56652 6072 56885 6100
rect 56652 6060 56658 6072
rect 56873 6069 56885 6072
rect 56919 6100 56931 6103
rect 57330 6100 57336 6112
rect 56919 6072 57336 6100
rect 56919 6069 56931 6072
rect 56873 6063 56931 6069
rect 57330 6060 57336 6072
rect 57388 6060 57394 6112
rect 57974 6100 57980 6112
rect 57935 6072 57980 6100
rect 57974 6060 57980 6072
rect 58032 6060 58038 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1854 5896 1860 5908
rect 1815 5868 1860 5896
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 56318 5760 56324 5772
rect 56279 5732 56324 5760
rect 56318 5720 56324 5732
rect 56376 5720 56382 5772
rect 56505 5763 56563 5769
rect 56505 5729 56517 5763
rect 56551 5760 56563 5763
rect 57974 5760 57980 5772
rect 56551 5732 57980 5760
rect 56551 5729 56563 5732
rect 56505 5723 56563 5729
rect 57974 5720 57980 5732
rect 58032 5720 58038 5772
rect 58158 5760 58164 5772
rect 58119 5732 58164 5760
rect 58158 5720 58164 5732
rect 58216 5720 58222 5772
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2096 5664 2329 5692
rect 2096 5652 2102 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2317 5655 2375 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 55490 5652 55496 5704
rect 55548 5692 55554 5704
rect 55861 5695 55919 5701
rect 55861 5692 55873 5695
rect 55548 5664 55873 5692
rect 55548 5652 55554 5664
rect 55861 5661 55873 5664
rect 55907 5661 55919 5695
rect 55861 5655 55919 5661
rect 3050 5556 3056 5568
rect 3011 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 3050 5284 3056 5296
rect 2179 5256 3056 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 55677 5287 55735 5293
rect 55677 5253 55689 5287
rect 55723 5284 55735 5287
rect 57054 5284 57060 5296
rect 55723 5256 57060 5284
rect 55723 5253 55735 5256
rect 55677 5247 55735 5253
rect 57054 5244 57060 5256
rect 57112 5244 57118 5296
rect 55490 5216 55496 5228
rect 55451 5188 55496 5216
rect 55490 5176 55496 5188
rect 55548 5176 55554 5228
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 1949 5151 2007 5157
rect 1949 5148 1961 5151
rect 1912 5120 1961 5148
rect 1912 5108 1918 5120
rect 1949 5117 1961 5120
rect 1995 5117 2007 5151
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 1949 5111 2007 5117
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 57333 5151 57391 5157
rect 57333 5117 57345 5151
rect 57379 5148 57391 5151
rect 58618 5148 58624 5160
rect 57379 5120 58624 5148
rect 57379 5117 57391 5120
rect 57333 5111 57391 5117
rect 58618 5108 58624 5120
rect 58676 5108 58682 5160
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 56318 4972 56324 5024
rect 56376 5012 56382 5024
rect 58069 5015 58127 5021
rect 58069 5012 58081 5015
rect 56376 4984 58081 5012
rect 56376 4972 56382 4984
rect 58069 4981 58081 4984
rect 58115 4981 58127 5015
rect 58069 4975 58127 4981
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1854 4808 1860 4820
rect 1815 4780 1860 4808
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 56318 4672 56324 4684
rect 56279 4644 56324 4672
rect 56318 4632 56324 4644
rect 56376 4632 56382 4684
rect 56502 4632 56508 4684
rect 56560 4672 56566 4684
rect 56781 4675 56839 4681
rect 56781 4672 56793 4675
rect 56560 4644 56793 4672
rect 56560 4632 56566 4644
rect 56781 4641 56793 4644
rect 56827 4641 56839 4675
rect 56781 4635 56839 4641
rect 2222 4564 2228 4616
rect 2280 4604 2286 4616
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2280 4576 2513 4604
rect 2280 4564 2286 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 7834 4604 7840 4616
rect 7795 4576 7840 4604
rect 2501 4567 2559 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 9122 4604 9128 4616
rect 9035 4576 9128 4604
rect 9122 4564 9128 4576
rect 9180 4604 9186 4616
rect 22830 4604 22836 4616
rect 9180 4576 22836 4604
rect 9180 4564 9186 4576
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 54757 4607 54815 4613
rect 54757 4573 54769 4607
rect 54803 4604 54815 4607
rect 55030 4604 55036 4616
rect 54803 4576 55036 4604
rect 54803 4573 54815 4576
rect 54757 4567 54815 4573
rect 55030 4564 55036 4576
rect 55088 4564 55094 4616
rect 55490 4564 55496 4616
rect 55548 4604 55554 4616
rect 55861 4607 55919 4613
rect 55861 4604 55873 4607
rect 55548 4576 55873 4604
rect 55548 4564 55554 4576
rect 55861 4573 55873 4576
rect 55907 4573 55919 4607
rect 55861 4567 55919 4573
rect 56505 4539 56563 4545
rect 56505 4505 56517 4539
rect 56551 4536 56563 4539
rect 57974 4536 57980 4548
rect 56551 4508 57980 4536
rect 56551 4505 56563 4508
rect 56505 4499 56563 4505
rect 57974 4496 57980 4508
rect 58032 4496 58038 4548
rect 7929 4471 7987 4477
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8202 4468 8208 4480
rect 7975 4440 8208 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 9217 4471 9275 4477
rect 9217 4437 9229 4471
rect 9263 4468 9275 4471
rect 9582 4468 9588 4480
rect 9263 4440 9588 4468
rect 9263 4437 9275 4440
rect 9217 4431 9275 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 8202 4196 8208 4208
rect 8163 4168 8208 4196
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 56594 4196 56600 4208
rect 30944 4168 31248 4196
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 14826 4128 14832 4140
rect 14787 4100 14832 4128
rect 7377 4091 7435 4097
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 1912 4032 2421 4060
rect 1912 4020 1918 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2774 4060 2780 4072
rect 2735 4032 2780 4060
rect 2409 4023 2467 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 7392 3992 7420 4091
rect 14826 4088 14832 4100
rect 14884 4128 14890 4140
rect 22462 4128 22468 4140
rect 14884 4100 16574 4128
rect 22423 4100 22468 4128
rect 14884 4088 14890 4100
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8294 4060 8300 4072
rect 8067 4032 8300 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8444 4032 8493 4060
rect 8444 4020 8450 4032
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 16546 4060 16574 4100
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 26970 4128 26976 4140
rect 26931 4100 26976 4128
rect 26970 4088 26976 4100
rect 27028 4088 27034 4140
rect 29822 4088 29828 4140
rect 29880 4128 29886 4140
rect 30944 4128 30972 4168
rect 31110 4128 31116 4140
rect 29880 4100 30972 4128
rect 31023 4100 31116 4128
rect 29880 4088 29886 4100
rect 31110 4088 31116 4100
rect 31168 4088 31174 4140
rect 31220 4128 31248 4168
rect 54772 4168 54984 4196
rect 38013 4131 38071 4137
rect 38013 4128 38025 4131
rect 31220 4100 38025 4128
rect 38013 4097 38025 4100
rect 38059 4097 38071 4131
rect 49970 4128 49976 4140
rect 38013 4091 38071 4097
rect 41386 4100 49976 4128
rect 29178 4060 29184 4072
rect 16546 4032 29184 4060
rect 8481 4023 8539 4029
rect 29178 4020 29184 4032
rect 29236 4020 29242 4072
rect 31128 4060 31156 4088
rect 31128 4032 35894 4060
rect 30558 3992 30564 4004
rect 7392 3964 30564 3992
rect 30558 3952 30564 3964
rect 30616 3952 30622 4004
rect 35866 3992 35894 4032
rect 41386 3992 41414 4100
rect 49970 4088 49976 4100
rect 50028 4088 50034 4140
rect 53834 4128 53840 4140
rect 53795 4100 53840 4128
rect 53834 4088 53840 4100
rect 53892 4128 53898 4140
rect 54772 4128 54800 4168
rect 53892 4100 54800 4128
rect 54849 4131 54907 4137
rect 53892 4088 53898 4100
rect 54849 4097 54861 4131
rect 54895 4097 54907 4131
rect 54956 4128 54984 4168
rect 55324 4168 56600 4196
rect 55324 4128 55352 4168
rect 56594 4156 56600 4168
rect 56652 4156 56658 4208
rect 55490 4128 55496 4140
rect 54956 4100 55352 4128
rect 55451 4100 55496 4128
rect 54849 4091 54907 4097
rect 46750 4020 46756 4072
rect 46808 4060 46814 4072
rect 54864 4060 54892 4091
rect 55490 4088 55496 4100
rect 55548 4088 55554 4140
rect 57790 4088 57796 4140
rect 57848 4128 57854 4140
rect 57885 4131 57943 4137
rect 57885 4128 57897 4131
rect 57848 4100 57897 4128
rect 57848 4088 57854 4100
rect 57885 4097 57897 4100
rect 57931 4097 57943 4131
rect 57885 4091 57943 4097
rect 46808 4032 54892 4060
rect 55691 4063 55749 4069
rect 46808 4020 46814 4032
rect 55691 4029 55703 4063
rect 55737 4029 55749 4063
rect 55691 4023 55749 4029
rect 57333 4063 57391 4069
rect 57333 4029 57345 4063
rect 57379 4060 57391 4063
rect 57698 4060 57704 4072
rect 57379 4032 57704 4060
rect 57379 4029 57391 4032
rect 57333 4023 57391 4029
rect 35866 3964 41414 3992
rect 44542 3952 44548 4004
rect 44600 3992 44606 4004
rect 55692 3992 55720 4023
rect 57698 4020 57704 4032
rect 57756 4020 57762 4072
rect 57977 3995 58035 4001
rect 57977 3992 57989 3995
rect 44600 3964 55628 3992
rect 55692 3964 57989 3992
rect 44600 3952 44606 3964
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 3844 3896 4721 3924
rect 3844 3884 3850 3896
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 7466 3924 7472 3936
rect 7427 3896 7472 3924
rect 4709 3887 4767 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 14921 3927 14979 3933
rect 14921 3893 14933 3927
rect 14967 3924 14979 3927
rect 15286 3924 15292 3936
rect 14967 3896 15292 3924
rect 14967 3893 14979 3896
rect 14921 3887 14979 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16853 3927 16911 3933
rect 16853 3924 16865 3927
rect 16724 3896 16865 3924
rect 16724 3884 16730 3896
rect 16853 3893 16865 3896
rect 16899 3893 16911 3927
rect 16853 3887 16911 3893
rect 22557 3927 22615 3933
rect 22557 3893 22569 3927
rect 22603 3924 22615 3927
rect 23014 3924 23020 3936
rect 22603 3896 23020 3924
rect 22603 3893 22615 3896
rect 22557 3887 22615 3893
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23290 3924 23296 3936
rect 23251 3896 23296 3924
rect 23290 3884 23296 3896
rect 23348 3884 23354 3936
rect 26878 3884 26884 3936
rect 26936 3924 26942 3936
rect 27065 3927 27123 3933
rect 27065 3924 27077 3927
rect 26936 3896 27077 3924
rect 26936 3884 26942 3896
rect 27065 3893 27077 3896
rect 27111 3893 27123 3927
rect 27065 3887 27123 3893
rect 29730 3884 29736 3936
rect 29788 3924 29794 3936
rect 30009 3927 30067 3933
rect 30009 3924 30021 3927
rect 29788 3896 30021 3924
rect 29788 3884 29794 3896
rect 30009 3893 30021 3896
rect 30055 3893 30067 3927
rect 30650 3924 30656 3936
rect 30611 3896 30656 3924
rect 30009 3887 30067 3893
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 30742 3884 30748 3936
rect 30800 3924 30806 3936
rect 31205 3927 31263 3933
rect 31205 3924 31217 3927
rect 30800 3896 31217 3924
rect 30800 3884 30806 3896
rect 31205 3893 31217 3896
rect 31251 3893 31263 3927
rect 31205 3887 31263 3893
rect 32122 3884 32128 3936
rect 32180 3924 32186 3936
rect 32309 3927 32367 3933
rect 32309 3924 32321 3927
rect 32180 3896 32321 3924
rect 32180 3884 32186 3896
rect 32309 3893 32321 3896
rect 32355 3893 32367 3927
rect 32309 3887 32367 3893
rect 38105 3927 38163 3933
rect 38105 3893 38117 3927
rect 38151 3924 38163 3927
rect 38470 3924 38476 3936
rect 38151 3896 38476 3924
rect 38151 3893 38163 3896
rect 38105 3887 38163 3893
rect 38470 3884 38476 3896
rect 38528 3884 38534 3936
rect 46290 3884 46296 3936
rect 46348 3924 46354 3936
rect 46477 3927 46535 3933
rect 46477 3924 46489 3927
rect 46348 3896 46489 3924
rect 46348 3884 46354 3896
rect 46477 3893 46489 3896
rect 46523 3893 46535 3927
rect 46477 3887 46535 3893
rect 50065 3927 50123 3933
rect 50065 3893 50077 3927
rect 50111 3924 50123 3927
rect 50338 3924 50344 3936
rect 50111 3896 50344 3924
rect 50111 3893 50123 3896
rect 50065 3887 50123 3893
rect 50338 3884 50344 3896
rect 50396 3884 50402 3936
rect 53098 3884 53104 3936
rect 53156 3924 53162 3936
rect 53929 3927 53987 3933
rect 53929 3924 53941 3927
rect 53156 3896 53941 3924
rect 53156 3884 53162 3896
rect 53929 3893 53941 3896
rect 53975 3893 53987 3927
rect 53929 3887 53987 3893
rect 54941 3927 54999 3933
rect 54941 3893 54953 3927
rect 54987 3924 54999 3927
rect 55398 3924 55404 3936
rect 54987 3896 55404 3924
rect 54987 3893 54999 3896
rect 54941 3887 54999 3893
rect 55398 3884 55404 3896
rect 55456 3884 55462 3936
rect 55600 3924 55628 3964
rect 57977 3961 57989 3964
rect 58023 3961 58035 3995
rect 57977 3955 58035 3961
rect 57146 3924 57152 3936
rect 55600 3896 57152 3924
rect 57146 3884 57152 3896
rect 57204 3884 57210 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 1854 3720 1860 3732
rect 1815 3692 1860 3720
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 8996 3692 16574 3720
rect 8996 3680 9002 3692
rect 16546 3652 16574 3692
rect 22462 3680 22468 3732
rect 22520 3720 22526 3732
rect 56778 3720 56784 3732
rect 22520 3692 56784 3720
rect 22520 3680 22526 3692
rect 56778 3680 56784 3692
rect 56836 3680 56842 3732
rect 22480 3652 22508 3680
rect 1780 3624 15424 3652
rect 16546 3624 22508 3652
rect 1780 3525 1808 3624
rect 3786 3584 3792 3596
rect 3747 3556 3792 3584
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4028 3556 4261 3584
rect 4028 3544 4034 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 5224 3556 6561 3584
rect 5224 3544 5230 3556
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 9582 3584 9588 3596
rect 9543 3556 9588 3584
rect 6549 3547 6607 3553
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9732 3556 9873 3584
rect 9732 3544 9738 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 15286 3584 15292 3596
rect 15247 3556 15292 3584
rect 9861 3547 9919 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15396 3584 15424 3624
rect 15396 3556 19656 3584
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2455 3488 3065 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 2314 3340 2320 3392
rect 2372 3380 2378 3392
rect 2501 3383 2559 3389
rect 2501 3380 2513 3383
rect 2372 3352 2513 3380
rect 2372 3340 2378 3352
rect 2501 3349 2513 3352
rect 2547 3349 2559 3383
rect 3068 3380 3096 3479
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5408 3488 6101 3516
rect 5408 3476 5414 3488
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3485 9459 3519
rect 12250 3516 12256 3528
rect 12211 3488 12256 3516
rect 9401 3479 9459 3485
rect 3145 3451 3203 3457
rect 3145 3417 3157 3451
rect 3191 3448 3203 3451
rect 3973 3451 4031 3457
rect 3973 3448 3985 3451
rect 3191 3420 3985 3448
rect 3191 3417 3203 3420
rect 3145 3411 3203 3417
rect 3973 3417 3985 3420
rect 4019 3417 4031 3451
rect 6270 3448 6276 3460
rect 6231 3420 6276 3448
rect 3973 3411 4031 3417
rect 6270 3408 6276 3420
rect 6328 3408 6334 3460
rect 9416 3448 9444 3479
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 12584 3488 13093 3516
rect 12584 3476 12590 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 15102 3516 15108 3528
rect 15063 3488 15108 3516
rect 13081 3479 13139 3485
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 17402 3516 17408 3528
rect 17363 3488 17408 3516
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 9766 3448 9772 3460
rect 9416 3420 9772 3448
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 15470 3408 15476 3460
rect 15528 3448 15534 3460
rect 16945 3451 17003 3457
rect 16945 3448 16957 3451
rect 15528 3420 16957 3448
rect 15528 3408 15534 3420
rect 16945 3417 16957 3420
rect 16991 3417 17003 3451
rect 16945 3411 17003 3417
rect 9214 3380 9220 3392
rect 3068 3352 9220 3380
rect 2501 3343 2559 3349
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 12345 3383 12403 3389
rect 12345 3349 12357 3383
rect 12391 3380 12403 3383
rect 12710 3380 12716 3392
rect 12391 3352 12716 3380
rect 12391 3349 12403 3352
rect 12345 3343 12403 3349
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 16850 3340 16856 3392
rect 16908 3380 16914 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 16908 3352 17509 3380
rect 16908 3340 16914 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 19628 3380 19656 3556
rect 19720 3525 19748 3624
rect 32950 3612 32956 3664
rect 33008 3652 33014 3664
rect 43254 3652 43260 3664
rect 33008 3624 43260 3652
rect 33008 3612 33014 3624
rect 43254 3612 43260 3624
rect 43312 3612 43318 3664
rect 57606 3652 57612 3664
rect 43456 3624 55214 3652
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20680 3556 20821 3584
rect 20680 3544 20686 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 25130 3584 25136 3596
rect 25091 3556 25136 3584
rect 20809 3547 20867 3553
rect 25130 3544 25136 3556
rect 25188 3544 25194 3596
rect 26878 3584 26884 3596
rect 26839 3556 26884 3584
rect 26878 3544 26884 3556
rect 26936 3544 26942 3596
rect 27062 3544 27068 3596
rect 27120 3584 27126 3596
rect 27157 3587 27215 3593
rect 27157 3584 27169 3587
rect 27120 3556 27169 3584
rect 27120 3544 27126 3556
rect 27157 3553 27169 3556
rect 27203 3553 27215 3587
rect 27157 3547 27215 3553
rect 29825 3587 29883 3593
rect 29825 3553 29837 3587
rect 29871 3584 29883 3587
rect 30650 3584 30656 3596
rect 29871 3556 30656 3584
rect 29871 3553 29883 3556
rect 29825 3547 29883 3553
rect 30650 3544 30656 3556
rect 30708 3544 30714 3596
rect 32122 3584 32128 3596
rect 32083 3556 32128 3584
rect 32122 3544 32128 3556
rect 32180 3544 32186 3596
rect 32858 3584 32864 3596
rect 32819 3556 32864 3584
rect 32858 3544 32864 3556
rect 32916 3544 32922 3596
rect 34146 3544 34152 3596
rect 34204 3584 34210 3596
rect 34204 3556 41276 3584
rect 34204 3544 34210 3556
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3485 19763 3519
rect 20346 3516 20352 3528
rect 20307 3488 20352 3516
rect 19705 3479 19763 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 22830 3516 22836 3528
rect 22791 3488 22836 3516
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 23891 3488 24409 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 26694 3516 26700 3528
rect 26655 3488 26700 3516
rect 24397 3479 24455 3485
rect 26694 3476 26700 3488
rect 26752 3476 26758 3528
rect 38286 3476 38292 3528
rect 38344 3516 38350 3528
rect 38565 3519 38623 3525
rect 38565 3516 38577 3519
rect 38344 3488 38577 3516
rect 38344 3476 38350 3488
rect 38565 3485 38577 3488
rect 38611 3485 38623 3519
rect 41248 3516 41276 3556
rect 43456 3516 43484 3624
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 47026 3584 47032 3596
rect 46987 3556 47032 3584
rect 47026 3544 47032 3556
rect 47084 3544 47090 3596
rect 50338 3584 50344 3596
rect 50299 3556 50344 3584
rect 50338 3544 50344 3556
rect 50396 3544 50402 3596
rect 50614 3584 50620 3596
rect 50575 3556 50620 3584
rect 50614 3544 50620 3556
rect 50672 3544 50678 3596
rect 53098 3584 53104 3596
rect 53059 3556 53104 3584
rect 53098 3544 53104 3556
rect 53156 3544 53162 3596
rect 54110 3584 54116 3596
rect 54071 3556 54116 3584
rect 54110 3544 54116 3556
rect 54168 3544 54174 3596
rect 41248 3488 43484 3516
rect 38565 3479 38623 3485
rect 48222 3476 48228 3528
rect 48280 3516 48286 3528
rect 48777 3519 48835 3525
rect 48777 3516 48789 3519
rect 48280 3488 48789 3516
rect 48280 3476 48286 3488
rect 48777 3485 48789 3488
rect 48823 3485 48835 3519
rect 48777 3479 48835 3485
rect 49605 3519 49663 3525
rect 49605 3485 49617 3519
rect 49651 3516 49663 3519
rect 50157 3519 50215 3525
rect 50157 3516 50169 3519
rect 49651 3488 50169 3516
rect 49651 3485 49663 3488
rect 49605 3479 49663 3485
rect 50157 3485 50169 3488
rect 50203 3485 50215 3519
rect 52914 3516 52920 3528
rect 52875 3488 52920 3516
rect 50157 3479 50215 3485
rect 52914 3476 52920 3488
rect 52972 3476 52978 3528
rect 19797 3451 19855 3457
rect 19797 3417 19809 3451
rect 19843 3448 19855 3451
rect 20533 3451 20591 3457
rect 20533 3448 20545 3451
rect 19843 3420 20545 3448
rect 19843 3417 19855 3420
rect 19797 3411 19855 3417
rect 20533 3417 20545 3420
rect 20579 3417 20591 3451
rect 20533 3411 20591 3417
rect 22925 3451 22983 3457
rect 22925 3417 22937 3451
rect 22971 3448 22983 3451
rect 24581 3451 24639 3457
rect 24581 3448 24593 3451
rect 22971 3420 24593 3448
rect 22971 3417 22983 3420
rect 22925 3411 22983 3417
rect 24581 3417 24593 3420
rect 24627 3417 24639 3451
rect 28810 3448 28816 3460
rect 24581 3411 24639 3417
rect 26206 3420 28816 3448
rect 26206 3380 26234 3420
rect 28810 3408 28816 3420
rect 28868 3408 28874 3460
rect 30009 3451 30067 3457
rect 30009 3417 30021 3451
rect 30055 3448 30067 3451
rect 31202 3448 31208 3460
rect 30055 3420 31208 3448
rect 30055 3417 30067 3420
rect 30009 3411 30067 3417
rect 31202 3408 31208 3420
rect 31260 3408 31266 3460
rect 31570 3408 31576 3460
rect 31628 3448 31634 3460
rect 31665 3451 31723 3457
rect 31665 3448 31677 3451
rect 31628 3420 31677 3448
rect 31628 3408 31634 3420
rect 31665 3417 31677 3420
rect 31711 3417 31723 3451
rect 31665 3411 31723 3417
rect 32309 3451 32367 3457
rect 32309 3417 32321 3451
rect 32355 3448 32367 3451
rect 32674 3448 32680 3460
rect 32355 3420 32680 3448
rect 32355 3417 32367 3420
rect 32309 3411 32367 3417
rect 32674 3408 32680 3420
rect 32732 3408 32738 3460
rect 43254 3408 43260 3460
rect 43312 3448 43318 3460
rect 46477 3451 46535 3457
rect 43312 3420 44680 3448
rect 43312 3408 43318 3420
rect 19628 3352 26234 3380
rect 17497 3343 17555 3349
rect 26970 3340 26976 3392
rect 27028 3380 27034 3392
rect 44542 3380 44548 3392
rect 27028 3352 44548 3380
rect 27028 3340 27034 3352
rect 44542 3340 44548 3352
rect 44600 3340 44606 3392
rect 44652 3380 44680 3420
rect 46477 3417 46489 3451
rect 46523 3448 46535 3451
rect 46842 3448 46848 3460
rect 46523 3420 46848 3448
rect 46523 3417 46535 3420
rect 46477 3411 46535 3417
rect 46842 3408 46848 3420
rect 46900 3408 46906 3460
rect 55186 3448 55214 3624
rect 55324 3624 57612 3652
rect 55324 3525 55352 3624
rect 57606 3612 57612 3624
rect 57664 3612 57670 3664
rect 56321 3587 56379 3593
rect 56321 3553 56333 3587
rect 56367 3584 56379 3587
rect 57882 3584 57888 3596
rect 56367 3556 57744 3584
rect 57843 3556 57888 3584
rect 56367 3553 56379 3556
rect 56321 3547 56379 3553
rect 55309 3519 55367 3525
rect 55309 3485 55321 3519
rect 55355 3485 55367 3519
rect 57716 3516 57744 3556
rect 57882 3544 57888 3556
rect 57940 3544 57946 3596
rect 58066 3516 58072 3528
rect 57716 3488 58072 3516
rect 55309 3479 55367 3485
rect 58066 3476 58072 3488
rect 58124 3476 58130 3528
rect 56042 3448 56048 3460
rect 55186 3420 56048 3448
rect 56042 3408 56048 3420
rect 56100 3408 56106 3460
rect 56505 3451 56563 3457
rect 56505 3417 56517 3451
rect 56551 3448 56563 3451
rect 56962 3448 56968 3460
rect 56551 3420 56968 3448
rect 56551 3417 56563 3420
rect 56505 3411 56563 3417
rect 56962 3408 56968 3420
rect 57020 3408 57026 3460
rect 48314 3380 48320 3392
rect 44652 3352 48320 3380
rect 48314 3340 48320 3352
rect 48372 3340 48378 3392
rect 54202 3340 54208 3392
rect 54260 3380 54266 3392
rect 55401 3383 55459 3389
rect 55401 3380 55413 3383
rect 54260 3352 55413 3380
rect 54260 3340 54266 3352
rect 55401 3349 55413 3352
rect 55447 3349 55459 3383
rect 55401 3343 55459 3349
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 6270 3176 6276 3188
rect 4663 3148 6276 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 23290 3176 23296 3188
rect 22848 3148 23296 3176
rect 2314 3108 2320 3120
rect 2275 3080 2320 3108
rect 2314 3068 2320 3080
rect 2372 3068 2378 3120
rect 12250 3108 12256 3120
rect 4724 3080 12256 3108
rect 4724 3052 4752 3080
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 12710 3108 12716 3120
rect 12671 3080 12716 3108
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 16850 3108 16856 3120
rect 16811 3080 16856 3108
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4706 3040 4712 3052
rect 4571 3012 4712 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5350 3040 5356 3052
rect 5311 3012 5356 3040
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 12526 3040 12532 3052
rect 12487 3012 12532 3040
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 15102 3000 15108 3052
rect 15160 3040 15166 3052
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 15160 3012 15393 3040
rect 15160 3000 15166 3012
rect 15381 3009 15393 3012
rect 15427 3009 15439 3043
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 15381 3003 15439 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 20346 3000 20352 3052
rect 20404 3040 20410 3052
rect 22848 3049 22876 3148
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 32674 3176 32680 3188
rect 32635 3148 32680 3176
rect 32674 3136 32680 3148
rect 32732 3136 32738 3188
rect 46842 3176 46848 3188
rect 46803 3148 46848 3176
rect 46842 3136 46848 3148
rect 46900 3136 46906 3188
rect 49970 3136 49976 3188
rect 50028 3176 50034 3188
rect 56962 3176 56968 3188
rect 50028 3148 55214 3176
rect 56923 3148 56968 3176
rect 50028 3136 50034 3148
rect 23014 3108 23020 3120
rect 22975 3080 23020 3108
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 29917 3111 29975 3117
rect 29917 3077 29929 3111
rect 29963 3108 29975 3111
rect 30742 3108 30748 3120
rect 29963 3080 30748 3108
rect 29963 3077 29975 3080
rect 29917 3071 29975 3077
rect 30742 3068 30748 3080
rect 30800 3068 30806 3120
rect 38470 3108 38476 3120
rect 38431 3080 38476 3108
rect 38470 3068 38476 3080
rect 38528 3068 38534 3120
rect 47673 3111 47731 3117
rect 47673 3077 47685 3111
rect 47719 3108 47731 3111
rect 48409 3111 48467 3117
rect 48409 3108 48421 3111
rect 47719 3080 48421 3108
rect 47719 3077 47731 3080
rect 47673 3071 47731 3077
rect 48409 3077 48421 3080
rect 48455 3077 48467 3111
rect 54202 3108 54208 3120
rect 54163 3080 54208 3108
rect 48409 3071 48467 3077
rect 54202 3068 54208 3080
rect 54260 3068 54266 3120
rect 55186 3108 55214 3148
rect 56962 3136 56968 3148
rect 57020 3136 57026 3188
rect 57974 3176 57980 3188
rect 57935 3148 57980 3176
rect 57974 3136 57980 3148
rect 58032 3136 58038 3188
rect 55186 3080 57928 3108
rect 20533 3043 20591 3049
rect 20533 3040 20545 3043
rect 20404 3012 20545 3040
rect 20404 3000 20410 3012
rect 20533 3009 20545 3012
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 26694 3000 26700 3052
rect 26752 3040 26758 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26752 3012 27169 3040
rect 26752 3000 26758 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 29730 3040 29736 3052
rect 29691 3012 29736 3040
rect 27157 3003 27215 3009
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 32585 3043 32643 3049
rect 32585 3040 32597 3043
rect 31128 3012 32597 3040
rect 2130 2972 2136 2984
rect 2091 2944 2136 2972
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2941 2651 2975
rect 2593 2935 2651 2941
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7607 2944 8033 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 8205 2975 8263 2981
rect 8205 2941 8217 2975
rect 8251 2972 8263 2975
rect 9030 2972 9036 2984
rect 8251 2944 9036 2972
rect 8251 2941 8263 2944
rect 8205 2935 8263 2941
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 2608 2904 2636 2935
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 716 2876 2636 2904
rect 716 2864 722 2876
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 9140 2904 9168 2935
rect 12894 2932 12900 2984
rect 12952 2972 12958 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12952 2944 13001 2972
rect 12952 2932 12958 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 16172 2944 17141 2972
rect 16172 2932 16178 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 23198 2932 23204 2984
rect 23256 2972 23262 2984
rect 23293 2975 23351 2981
rect 23293 2972 23305 2975
rect 23256 2944 23305 2972
rect 23256 2932 23262 2944
rect 23293 2941 23305 2944
rect 23339 2941 23351 2975
rect 30926 2972 30932 2984
rect 30887 2944 30932 2972
rect 23293 2935 23351 2941
rect 30926 2932 30932 2944
rect 30984 2932 30990 2984
rect 7800 2876 9168 2904
rect 7800 2864 7806 2876
rect 31128 2848 31156 3012
rect 32585 3009 32597 3012
rect 32631 3009 32643 3043
rect 38286 3040 38292 3052
rect 38247 3012 38292 3040
rect 32585 3003 32643 3009
rect 38286 3000 38292 3012
rect 38344 3000 38350 3052
rect 46750 3040 46756 3052
rect 46711 3012 46756 3040
rect 46750 3000 46756 3012
rect 46808 3000 46814 3052
rect 47578 3040 47584 3052
rect 47539 3012 47584 3040
rect 47578 3000 47584 3012
rect 47636 3000 47642 3052
rect 48222 3040 48228 3052
rect 48183 3012 48228 3040
rect 48222 3000 48228 3012
rect 48280 3000 48286 3052
rect 52914 3000 52920 3052
rect 52972 3040 52978 3052
rect 53561 3043 53619 3049
rect 53561 3040 53573 3043
rect 52972 3012 53573 3040
rect 52972 3000 52978 3012
rect 53561 3009 53573 3012
rect 53607 3009 53619 3043
rect 53561 3003 53619 3009
rect 56778 3000 56784 3052
rect 56836 3040 56842 3052
rect 57900 3049 57928 3080
rect 56873 3043 56931 3049
rect 56873 3040 56885 3043
rect 56836 3012 56885 3040
rect 56836 3000 56842 3012
rect 56873 3009 56885 3012
rect 56919 3009 56931 3043
rect 56873 3003 56931 3009
rect 57885 3043 57943 3049
rect 57885 3009 57897 3043
rect 57931 3009 57943 3043
rect 57885 3003 57943 3009
rect 38654 2932 38660 2984
rect 38712 2972 38718 2984
rect 38749 2975 38807 2981
rect 38749 2972 38761 2975
rect 38712 2944 38761 2972
rect 38712 2932 38718 2944
rect 38749 2941 38761 2944
rect 38795 2941 38807 2975
rect 49602 2972 49608 2984
rect 49563 2944 49608 2972
rect 38749 2935 38807 2941
rect 49602 2932 49608 2944
rect 49660 2932 49666 2984
rect 54018 2972 54024 2984
rect 53979 2944 54024 2972
rect 54018 2932 54024 2944
rect 54076 2932 54082 2984
rect 54754 2972 54760 2984
rect 54715 2944 54760 2972
rect 54754 2932 54760 2944
rect 54812 2932 54818 2984
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 6972 2808 7017 2836
rect 6972 2796 6978 2808
rect 28810 2796 28816 2848
rect 28868 2836 28874 2848
rect 31110 2836 31116 2848
rect 28868 2808 31116 2836
rect 28868 2796 28874 2808
rect 31110 2796 31116 2808
rect 31168 2796 31174 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2188 2604 2421 2632
rect 2188 2592 2194 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 9030 2632 9036 2644
rect 8991 2604 9036 2632
rect 2409 2595 2467 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 31202 2632 31208 2644
rect 31163 2604 31208 2632
rect 31202 2592 31208 2604
rect 31260 2592 31266 2644
rect 54018 2592 54024 2644
rect 54076 2632 54082 2644
rect 54205 2635 54263 2641
rect 54205 2632 54217 2635
rect 54076 2604 54217 2632
rect 54076 2592 54082 2604
rect 54205 2601 54217 2604
rect 54251 2601 54263 2635
rect 58066 2632 58072 2644
rect 58027 2604 58072 2632
rect 54205 2595 54263 2601
rect 58066 2592 58072 2604
rect 58124 2592 58130 2644
rect 6454 2524 6460 2576
rect 6512 2564 6518 2576
rect 6512 2536 7052 2564
rect 6512 2524 6518 2536
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 6914 2496 6920 2508
rect 6595 2468 6920 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7024 2505 7052 2536
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 53834 2496 53840 2508
rect 7009 2459 7067 2465
rect 16546 2468 53840 2496
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2428 8999 2431
rect 16546 2428 16574 2468
rect 53834 2456 53840 2468
rect 53892 2456 53898 2508
rect 55030 2456 55036 2508
rect 55088 2496 55094 2508
rect 55493 2499 55551 2505
rect 55493 2496 55505 2499
rect 55088 2468 55505 2496
rect 55088 2456 55094 2468
rect 55493 2465 55505 2468
rect 55539 2465 55551 2499
rect 55493 2459 55551 2465
rect 31110 2428 31116 2440
rect 8987 2400 16574 2428
rect 31071 2400 31116 2428
rect 8987 2397 8999 2400
rect 8941 2391 8999 2397
rect 31110 2388 31116 2400
rect 31168 2388 31174 2440
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7466 2360 7472 2372
rect 6779 2332 7472 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 55398 2320 55404 2372
rect 55456 2360 55462 2372
rect 55677 2363 55735 2369
rect 55677 2360 55689 2363
rect 55456 2332 55689 2360
rect 55456 2320 55462 2332
rect 55677 2329 55689 2332
rect 55723 2329 55735 2363
rect 57330 2360 57336 2372
rect 57291 2332 57336 2360
rect 55677 2323 55735 2329
rect 57330 2320 57336 2332
rect 57388 2320 57394 2372
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 664 57400 716 57452
rect 10324 57400 10376 57452
rect 33508 57400 33560 57452
rect 57704 57400 57756 57452
rect 20444 57332 20496 57384
rect 22008 57264 22060 57316
rect 3700 57196 3752 57248
rect 3792 57196 3844 57248
rect 17960 57239 18012 57248
rect 17960 57205 17969 57239
rect 17969 57205 18003 57239
rect 18003 57205 18012 57239
rect 17960 57196 18012 57205
rect 18052 57196 18104 57248
rect 19248 57196 19300 57248
rect 31300 57196 31352 57248
rect 32128 57196 32180 57248
rect 33600 57239 33652 57248
rect 33600 57205 33609 57239
rect 33609 57205 33643 57239
rect 33643 57205 33652 57239
rect 33600 57196 33652 57205
rect 35624 57196 35676 57248
rect 56324 57196 56376 57248
rect 56600 57196 56652 57248
rect 57244 57239 57296 57248
rect 57244 57205 57253 57239
rect 57253 57205 57287 57239
rect 57287 57205 57296 57239
rect 57244 57196 57296 57205
rect 57428 57196 57480 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 3792 56899 3844 56908
rect 3792 56865 3801 56899
rect 3801 56865 3835 56899
rect 3835 56865 3844 56899
rect 3792 56856 3844 56865
rect 4160 56856 4212 56908
rect 1952 56788 2004 56840
rect 2872 56831 2924 56840
rect 2872 56797 2881 56831
rect 2881 56797 2915 56831
rect 2915 56797 2924 56831
rect 2872 56788 2924 56797
rect 6368 56788 6420 56840
rect 8668 56788 8720 56840
rect 13268 56788 13320 56840
rect 16028 56831 16080 56840
rect 16028 56797 16037 56831
rect 16037 56797 16071 56831
rect 16071 56797 16080 56831
rect 16028 56788 16080 56797
rect 17316 56788 17368 56840
rect 46664 56856 46716 56908
rect 56324 56899 56376 56908
rect 56324 56865 56333 56899
rect 56333 56865 56367 56899
rect 56367 56865 56376 56899
rect 56324 56856 56376 56865
rect 57980 56899 58032 56908
rect 57980 56865 57989 56899
rect 57989 56865 58023 56899
rect 58023 56865 58032 56899
rect 57980 56856 58032 56865
rect 18236 56831 18288 56840
rect 18236 56797 18245 56831
rect 18245 56797 18279 56831
rect 18279 56797 18288 56831
rect 18236 56788 18288 56797
rect 22560 56831 22612 56840
rect 22560 56797 22569 56831
rect 22569 56797 22603 56831
rect 22603 56797 22612 56831
rect 22560 56788 22612 56797
rect 27252 56831 27304 56840
rect 27252 56797 27261 56831
rect 27261 56797 27295 56831
rect 27295 56797 27304 56831
rect 27252 56788 27304 56797
rect 27896 56831 27948 56840
rect 27896 56797 27905 56831
rect 27905 56797 27939 56831
rect 27939 56797 27948 56831
rect 27896 56788 27948 56797
rect 28264 56788 28316 56840
rect 30196 56831 30248 56840
rect 30196 56797 30205 56831
rect 30205 56797 30239 56831
rect 30239 56797 30248 56831
rect 30196 56788 30248 56797
rect 30656 56831 30708 56840
rect 30656 56797 30665 56831
rect 30665 56797 30699 56831
rect 30699 56797 30708 56831
rect 30656 56788 30708 56797
rect 31300 56831 31352 56840
rect 31300 56797 31309 56831
rect 31309 56797 31343 56831
rect 31343 56797 31352 56831
rect 31300 56788 31352 56797
rect 35624 56831 35676 56840
rect 35624 56797 35633 56831
rect 35633 56797 35667 56831
rect 35667 56797 35676 56831
rect 35624 56788 35676 56797
rect 40040 56831 40092 56840
rect 40040 56797 40049 56831
rect 40049 56797 40083 56831
rect 40083 56797 40092 56831
rect 40040 56788 40092 56797
rect 42248 56831 42300 56840
rect 42248 56797 42257 56831
rect 42257 56797 42291 56831
rect 42291 56797 42300 56831
rect 42248 56788 42300 56797
rect 42892 56831 42944 56840
rect 42892 56797 42901 56831
rect 42901 56797 42935 56831
rect 42935 56797 42944 56831
rect 42892 56788 42944 56797
rect 46204 56788 46256 56840
rect 49700 56788 49752 56840
rect 55496 56788 55548 56840
rect 4344 56720 4396 56772
rect 31760 56720 31812 56772
rect 35808 56763 35860 56772
rect 35808 56729 35817 56763
rect 35817 56729 35851 56763
rect 35851 56729 35860 56763
rect 35808 56720 35860 56729
rect 36084 56720 36136 56772
rect 57980 56720 58032 56772
rect 17868 56652 17920 56704
rect 22376 56695 22428 56704
rect 22376 56661 22385 56695
rect 22385 56661 22419 56695
rect 22419 56661 22428 56695
rect 22376 56652 22428 56661
rect 27160 56652 27212 56704
rect 28172 56652 28224 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4344 56491 4396 56500
rect 4344 56457 4353 56491
rect 4353 56457 4387 56491
rect 4387 56457 4396 56491
rect 4344 56448 4396 56457
rect 22560 56448 22612 56500
rect 26976 56448 27028 56500
rect 27252 56448 27304 56500
rect 1952 56355 2004 56364
rect 1952 56321 1961 56355
rect 1961 56321 1995 56355
rect 1995 56321 2004 56355
rect 1952 56312 2004 56321
rect 6368 56355 6420 56364
rect 2136 56287 2188 56296
rect 2136 56253 2145 56287
rect 2145 56253 2179 56287
rect 2179 56253 2188 56287
rect 2136 56244 2188 56253
rect 2780 56287 2832 56296
rect 2780 56253 2789 56287
rect 2789 56253 2823 56287
rect 2823 56253 2832 56287
rect 2780 56244 2832 56253
rect 6368 56321 6377 56355
rect 6377 56321 6411 56355
rect 6411 56321 6420 56355
rect 6368 56312 6420 56321
rect 8668 56355 8720 56364
rect 8668 56321 8677 56355
rect 8677 56321 8711 56355
rect 8711 56321 8720 56355
rect 8668 56312 8720 56321
rect 13268 56355 13320 56364
rect 13268 56321 13277 56355
rect 13277 56321 13311 56355
rect 13311 56321 13320 56355
rect 13268 56312 13320 56321
rect 18236 56380 18288 56432
rect 22376 56380 22428 56432
rect 28172 56423 28224 56432
rect 28172 56389 28181 56423
rect 28181 56389 28215 56423
rect 28215 56389 28224 56423
rect 28172 56380 28224 56389
rect 30656 56380 30708 56432
rect 22008 56355 22060 56364
rect 22008 56321 22017 56355
rect 22017 56321 22051 56355
rect 22051 56321 22060 56355
rect 22008 56312 22060 56321
rect 26148 56312 26200 56364
rect 27896 56312 27948 56364
rect 31484 56380 31536 56432
rect 47860 56448 47912 56500
rect 32128 56355 32180 56364
rect 32128 56321 32137 56355
rect 32137 56321 32171 56355
rect 32171 56321 32180 56355
rect 32128 56312 32180 56321
rect 40040 56380 40092 56432
rect 42892 56380 42944 56432
rect 44456 56423 44508 56432
rect 44456 56389 44465 56423
rect 44465 56389 44499 56423
rect 44499 56389 44508 56423
rect 44456 56380 44508 56389
rect 46664 56355 46716 56364
rect 46664 56321 46673 56355
rect 46673 56321 46707 56355
rect 46707 56321 46716 56355
rect 46664 56312 46716 56321
rect 49700 56380 49752 56432
rect 55496 56355 55548 56364
rect 55496 56321 55505 56355
rect 55505 56321 55539 56355
rect 55539 56321 55548 56355
rect 55496 56312 55548 56321
rect 56876 56312 56928 56364
rect 6920 56244 6972 56296
rect 5816 56176 5868 56228
rect 9036 56244 9088 56296
rect 7104 56176 7156 56228
rect 13084 56244 13136 56296
rect 13544 56244 13596 56296
rect 17132 56244 17184 56296
rect 17408 56287 17460 56296
rect 17408 56253 17417 56287
rect 17417 56253 17451 56287
rect 17451 56253 17460 56287
rect 17408 56244 17460 56253
rect 19064 56287 19116 56296
rect 19064 56253 19073 56287
rect 19073 56253 19107 56287
rect 19107 56253 19116 56287
rect 19064 56244 19116 56253
rect 4712 56108 4764 56160
rect 15108 56108 15160 56160
rect 19340 56244 19392 56296
rect 21824 56287 21876 56296
rect 21824 56253 21833 56287
rect 21833 56253 21867 56287
rect 21867 56253 21876 56287
rect 21824 56244 21876 56253
rect 23020 56287 23072 56296
rect 23020 56253 23029 56287
rect 23029 56253 23063 56287
rect 23063 56253 23072 56287
rect 23020 56244 23072 56253
rect 26976 56287 27028 56296
rect 26976 56253 26985 56287
rect 26985 56253 27019 56287
rect 27019 56253 27028 56287
rect 26976 56244 27028 56253
rect 28356 56244 28408 56296
rect 32404 56244 32456 56296
rect 32864 56287 32916 56296
rect 32864 56253 32873 56287
rect 32873 56253 32907 56287
rect 32907 56253 32916 56287
rect 32864 56244 32916 56253
rect 40132 56244 40184 56296
rect 40592 56287 40644 56296
rect 40592 56253 40601 56287
rect 40601 56253 40635 56287
rect 40635 56253 40644 56287
rect 40592 56244 40644 56253
rect 42800 56287 42852 56296
rect 42800 56253 42809 56287
rect 42809 56253 42843 56287
rect 42843 56253 42852 56287
rect 42800 56244 42852 56253
rect 50252 56244 50304 56296
rect 56692 56287 56744 56296
rect 27620 56176 27672 56228
rect 50160 56176 50212 56228
rect 56692 56253 56701 56287
rect 56701 56253 56735 56287
rect 56735 56253 56744 56287
rect 56692 56244 56744 56253
rect 19340 56108 19392 56160
rect 25596 56108 25648 56160
rect 30932 56151 30984 56160
rect 30932 56117 30941 56151
rect 30941 56117 30975 56151
rect 30975 56117 30984 56151
rect 30932 56108 30984 56117
rect 35716 56108 35768 56160
rect 46388 56108 46440 56160
rect 56232 56108 56284 56160
rect 56876 56108 56928 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 6920 55904 6972 55956
rect 9036 55947 9088 55956
rect 9036 55913 9045 55947
rect 9045 55913 9079 55947
rect 9079 55913 9088 55947
rect 9036 55904 9088 55913
rect 13084 55947 13136 55956
rect 13084 55913 13093 55947
rect 13093 55913 13127 55947
rect 13127 55913 13136 55947
rect 13084 55904 13136 55913
rect 50252 55947 50304 55956
rect 9496 55836 9548 55888
rect 19064 55836 19116 55888
rect 20444 55879 20496 55888
rect 20444 55845 20453 55879
rect 20453 55845 20487 55879
rect 20487 55845 20496 55879
rect 20444 55836 20496 55845
rect 28172 55836 28224 55888
rect 32404 55879 32456 55888
rect 1492 55743 1544 55752
rect 1492 55709 1501 55743
rect 1501 55709 1535 55743
rect 1535 55709 1544 55743
rect 1492 55700 1544 55709
rect 3700 55700 3752 55752
rect 2044 55675 2096 55684
rect 2044 55641 2053 55675
rect 2053 55641 2087 55675
rect 2087 55641 2096 55675
rect 2044 55632 2096 55641
rect 2596 55564 2648 55616
rect 16028 55768 16080 55820
rect 16120 55768 16172 55820
rect 8944 55743 8996 55752
rect 8944 55709 8953 55743
rect 8953 55709 8987 55743
rect 8987 55709 8996 55743
rect 8944 55700 8996 55709
rect 12992 55743 13044 55752
rect 12992 55709 13001 55743
rect 13001 55709 13035 55743
rect 13035 55709 13044 55743
rect 12992 55700 13044 55709
rect 15108 55743 15160 55752
rect 15108 55709 15117 55743
rect 15117 55709 15151 55743
rect 15151 55709 15160 55743
rect 15108 55700 15160 55709
rect 21824 55743 21876 55752
rect 21824 55709 21833 55743
rect 21833 55709 21867 55743
rect 21867 55709 21876 55743
rect 21824 55700 21876 55709
rect 16580 55564 16632 55616
rect 17316 55564 17368 55616
rect 21272 55564 21324 55616
rect 22560 55607 22612 55616
rect 22560 55573 22569 55607
rect 22569 55573 22603 55607
rect 22603 55573 22612 55607
rect 22560 55564 22612 55573
rect 23020 55768 23072 55820
rect 30196 55768 30248 55820
rect 30288 55768 30340 55820
rect 32404 55845 32413 55879
rect 32413 55845 32447 55879
rect 32447 55845 32456 55879
rect 32404 55836 32456 55845
rect 35808 55836 35860 55888
rect 40132 55879 40184 55888
rect 40132 55845 40141 55879
rect 40141 55845 40175 55879
rect 40175 55845 40184 55879
rect 40132 55836 40184 55845
rect 50252 55913 50261 55947
rect 50261 55913 50295 55947
rect 50295 55913 50304 55947
rect 50252 55904 50304 55913
rect 55404 55904 55456 55956
rect 57244 55904 57296 55956
rect 42248 55768 42300 55820
rect 43812 55811 43864 55820
rect 43812 55777 43821 55811
rect 43821 55777 43855 55811
rect 43855 55777 43864 55811
rect 43812 55768 43864 55777
rect 25044 55700 25096 55752
rect 27160 55700 27212 55752
rect 32220 55700 32272 55752
rect 35348 55700 35400 55752
rect 35716 55743 35768 55752
rect 35716 55709 35725 55743
rect 35725 55709 35759 55743
rect 35759 55709 35768 55743
rect 35716 55700 35768 55709
rect 40040 55743 40092 55752
rect 40040 55709 40049 55743
rect 40049 55709 40083 55743
rect 40083 55709 40092 55743
rect 40040 55700 40092 55709
rect 25412 55632 25464 55684
rect 26332 55607 26384 55616
rect 26332 55573 26341 55607
rect 26341 55573 26375 55607
rect 26375 55573 26384 55607
rect 26332 55564 26384 55573
rect 28448 55607 28500 55616
rect 28448 55573 28457 55607
rect 28457 55573 28491 55607
rect 28491 55573 28500 55607
rect 28448 55564 28500 55573
rect 30932 55632 30984 55684
rect 33600 55564 33652 55616
rect 36268 55632 36320 55684
rect 36728 55632 36780 55684
rect 42616 55675 42668 55684
rect 42616 55641 42625 55675
rect 42625 55641 42659 55675
rect 42659 55641 42668 55675
rect 42616 55632 42668 55641
rect 42800 55564 42852 55616
rect 56232 55836 56284 55888
rect 46204 55811 46256 55820
rect 46204 55777 46213 55811
rect 46213 55777 46247 55811
rect 46247 55777 46256 55811
rect 46204 55768 46256 55777
rect 46388 55811 46440 55820
rect 46388 55777 46397 55811
rect 46397 55777 46431 55811
rect 46431 55777 46440 55811
rect 46388 55768 46440 55777
rect 47032 55811 47084 55820
rect 47032 55777 47041 55811
rect 47041 55777 47075 55811
rect 47075 55777 47084 55811
rect 47032 55768 47084 55777
rect 56048 55768 56100 55820
rect 57428 55836 57480 55888
rect 56508 55768 56560 55820
rect 47860 55700 47912 55752
rect 52920 55743 52972 55752
rect 52920 55709 52929 55743
rect 52929 55709 52963 55743
rect 52963 55709 52972 55743
rect 52920 55700 52972 55709
rect 55312 55700 55364 55752
rect 55680 55743 55732 55752
rect 55680 55709 55689 55743
rect 55689 55709 55723 55743
rect 55723 55709 55732 55743
rect 55680 55700 55732 55709
rect 54668 55632 54720 55684
rect 56784 55564 56836 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 21824 55360 21876 55412
rect 2872 55292 2924 55344
rect 17960 55292 18012 55344
rect 22560 55292 22612 55344
rect 23664 55360 23716 55412
rect 25412 55403 25464 55412
rect 25412 55369 25421 55403
rect 25421 55369 25455 55403
rect 25455 55369 25464 55403
rect 25412 55360 25464 55369
rect 36268 55403 36320 55412
rect 27344 55292 27396 55344
rect 21272 55267 21324 55276
rect 21272 55233 21281 55267
rect 21281 55233 21315 55267
rect 21315 55233 21324 55267
rect 21272 55224 21324 55233
rect 21916 55224 21968 55276
rect 25596 55267 25648 55276
rect 25596 55233 25605 55267
rect 25605 55233 25639 55267
rect 25639 55233 25648 55267
rect 25596 55224 25648 55233
rect 26148 55224 26200 55276
rect 28540 55292 28592 55344
rect 29276 55224 29328 55276
rect 36268 55369 36277 55403
rect 36277 55369 36311 55403
rect 36311 55369 36320 55403
rect 36268 55360 36320 55369
rect 40040 55360 40092 55412
rect 54668 55403 54720 55412
rect 54668 55369 54677 55403
rect 54677 55369 54711 55403
rect 54711 55369 54720 55403
rect 54668 55360 54720 55369
rect 55312 55292 55364 55344
rect 36176 55267 36228 55276
rect 36176 55233 36185 55267
rect 36185 55233 36219 55267
rect 36219 55233 36228 55267
rect 36176 55224 36228 55233
rect 3792 55156 3844 55208
rect 3976 55199 4028 55208
rect 3976 55165 3985 55199
rect 3985 55165 4019 55199
rect 4019 55165 4028 55199
rect 3976 55156 4028 55165
rect 17868 55199 17920 55208
rect 17868 55165 17877 55199
rect 17877 55165 17911 55199
rect 17911 55165 17920 55199
rect 17868 55156 17920 55165
rect 19248 55199 19300 55208
rect 19248 55165 19257 55199
rect 19257 55165 19291 55199
rect 19291 55165 19300 55199
rect 19248 55156 19300 55165
rect 26056 55199 26108 55208
rect 26056 55165 26065 55199
rect 26065 55165 26099 55199
rect 26099 55165 26108 55199
rect 26056 55156 26108 55165
rect 28540 55156 28592 55208
rect 29552 55156 29604 55208
rect 29276 55131 29328 55140
rect 29276 55097 29285 55131
rect 29285 55097 29319 55131
rect 29319 55097 29328 55131
rect 29276 55088 29328 55097
rect 55404 55224 55456 55276
rect 56600 55360 56652 55412
rect 56784 55360 56836 55412
rect 57980 55403 58032 55412
rect 57336 55335 57388 55344
rect 57336 55301 57345 55335
rect 57345 55301 57379 55335
rect 57379 55301 57388 55335
rect 57336 55292 57388 55301
rect 57980 55369 57989 55403
rect 57989 55369 58023 55403
rect 58023 55369 58032 55403
rect 57980 55360 58032 55369
rect 56600 55088 56652 55140
rect 21088 55063 21140 55072
rect 21088 55029 21097 55063
rect 21097 55029 21131 55063
rect 21131 55029 21140 55063
rect 21088 55020 21140 55029
rect 27620 55020 27672 55072
rect 28080 55020 28132 55072
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 2136 54816 2188 54868
rect 3792 54816 3844 54868
rect 19340 54859 19392 54868
rect 19340 54825 19349 54859
rect 19349 54825 19383 54859
rect 19383 54825 19392 54859
rect 19340 54816 19392 54825
rect 27620 54816 27672 54868
rect 27896 54816 27948 54868
rect 28448 54816 28500 54868
rect 26056 54680 26108 54732
rect 29000 54680 29052 54732
rect 58164 54723 58216 54732
rect 58164 54689 58173 54723
rect 58173 54689 58207 54723
rect 58207 54689 58216 54723
rect 58164 54680 58216 54689
rect 3332 54612 3384 54664
rect 3976 54612 4028 54664
rect 19156 54612 19208 54664
rect 21916 54612 21968 54664
rect 21088 54544 21140 54596
rect 26976 54544 27028 54596
rect 29552 54655 29604 54664
rect 29552 54621 29561 54655
rect 29561 54621 29595 54655
rect 29595 54621 29604 54655
rect 29552 54612 29604 54621
rect 56324 54655 56376 54664
rect 56324 54621 56333 54655
rect 56333 54621 56367 54655
rect 56367 54621 56376 54655
rect 56324 54612 56376 54621
rect 28080 54587 28132 54596
rect 28080 54553 28089 54587
rect 28089 54553 28123 54587
rect 28123 54553 28132 54587
rect 28080 54544 28132 54553
rect 29644 54544 29696 54596
rect 34428 54544 34480 54596
rect 56968 54544 57020 54596
rect 19984 54476 20036 54528
rect 27436 54519 27488 54528
rect 27436 54485 27461 54519
rect 27461 54485 27488 54519
rect 27436 54476 27488 54485
rect 28448 54476 28500 54528
rect 28724 54476 28776 54528
rect 29000 54476 29052 54528
rect 52920 54476 52972 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 29644 54315 29696 54324
rect 29644 54281 29653 54315
rect 29653 54281 29687 54315
rect 29687 54281 29696 54315
rect 29644 54272 29696 54281
rect 56968 54315 57020 54324
rect 56968 54281 56977 54315
rect 56977 54281 57011 54315
rect 57011 54281 57020 54315
rect 56968 54272 57020 54281
rect 26332 54204 26384 54256
rect 26148 54136 26200 54188
rect 27896 54179 27948 54188
rect 27896 54145 27905 54179
rect 27905 54145 27939 54179
rect 27939 54145 27948 54179
rect 27896 54136 27948 54145
rect 29184 54204 29236 54256
rect 28448 54136 28500 54188
rect 56324 54204 56376 54256
rect 56232 54179 56284 54188
rect 29000 54111 29052 54120
rect 29000 54077 29009 54111
rect 29009 54077 29043 54111
rect 29043 54077 29052 54111
rect 29000 54068 29052 54077
rect 29092 54111 29144 54120
rect 29092 54077 29101 54111
rect 29101 54077 29135 54111
rect 29135 54077 29144 54111
rect 29092 54068 29144 54077
rect 56232 54145 56241 54179
rect 56241 54145 56275 54179
rect 56275 54145 56284 54179
rect 56232 54136 56284 54145
rect 56876 54179 56928 54188
rect 56876 54145 56885 54179
rect 56885 54145 56919 54179
rect 56919 54145 56928 54179
rect 56876 54136 56928 54145
rect 26240 53975 26292 53984
rect 26240 53941 26249 53975
rect 26249 53941 26283 53975
rect 26283 53941 26292 53975
rect 26240 53932 26292 53941
rect 29644 53932 29696 53984
rect 56508 53932 56560 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 27436 53728 27488 53780
rect 29092 53728 29144 53780
rect 26332 53660 26384 53712
rect 27252 53660 27304 53712
rect 25044 53592 25096 53644
rect 56508 53635 56560 53644
rect 56508 53601 56517 53635
rect 56517 53601 56551 53635
rect 56551 53601 56560 53635
rect 56508 53592 56560 53601
rect 58164 53635 58216 53644
rect 58164 53601 58173 53635
rect 58173 53601 58207 53635
rect 58207 53601 58216 53635
rect 58164 53592 58216 53601
rect 1952 53524 2004 53576
rect 22560 53567 22612 53576
rect 22560 53533 22569 53567
rect 22569 53533 22603 53567
rect 22603 53533 22612 53567
rect 22560 53524 22612 53533
rect 22744 53567 22796 53576
rect 22744 53533 22753 53567
rect 22753 53533 22787 53567
rect 22787 53533 22796 53567
rect 22744 53524 22796 53533
rect 26792 53524 26844 53576
rect 27436 53524 27488 53576
rect 28724 53567 28776 53576
rect 28724 53533 28733 53567
rect 28733 53533 28767 53567
rect 28767 53533 28776 53567
rect 28724 53524 28776 53533
rect 29000 53567 29052 53576
rect 25412 53499 25464 53508
rect 25412 53465 25446 53499
rect 25446 53465 25464 53499
rect 25412 53456 25464 53465
rect 26884 53456 26936 53508
rect 28448 53456 28500 53508
rect 29000 53533 29009 53567
rect 29009 53533 29043 53567
rect 29043 53533 29052 53567
rect 29000 53524 29052 53533
rect 29552 53567 29604 53576
rect 29552 53533 29561 53567
rect 29561 53533 29595 53567
rect 29595 53533 29604 53567
rect 29552 53524 29604 53533
rect 29644 53524 29696 53576
rect 56324 53567 56376 53576
rect 56324 53533 56333 53567
rect 56333 53533 56367 53567
rect 56367 53533 56376 53567
rect 56324 53524 56376 53533
rect 22376 53388 22428 53440
rect 27160 53431 27212 53440
rect 27160 53397 27169 53431
rect 27169 53397 27203 53431
rect 27203 53397 27212 53431
rect 27160 53388 27212 53397
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 25412 53227 25464 53236
rect 25412 53193 25421 53227
rect 25421 53193 25455 53227
rect 25455 53193 25464 53227
rect 25412 53184 25464 53193
rect 27436 53227 27488 53236
rect 5172 53116 5224 53168
rect 25780 53116 25832 53168
rect 27436 53193 27445 53227
rect 27445 53193 27479 53227
rect 27479 53193 27488 53227
rect 27436 53184 27488 53193
rect 1952 53091 2004 53100
rect 1952 53057 1961 53091
rect 1961 53057 1995 53091
rect 1995 53057 2004 53091
rect 1952 53048 2004 53057
rect 21916 53048 21968 53100
rect 22100 53091 22152 53100
rect 22100 53057 22134 53091
rect 22134 53057 22152 53091
rect 23664 53091 23716 53100
rect 22100 53048 22152 53057
rect 23664 53057 23673 53091
rect 23673 53057 23707 53091
rect 23707 53057 23716 53091
rect 23664 53048 23716 53057
rect 25504 53048 25556 53100
rect 26148 53048 26200 53100
rect 28172 53116 28224 53168
rect 26884 53048 26936 53100
rect 27252 53091 27304 53100
rect 27252 53057 27261 53091
rect 27261 53057 27295 53091
rect 27295 53057 27304 53091
rect 27252 53048 27304 53057
rect 27344 53048 27396 53100
rect 56324 53048 56376 53100
rect 2412 52980 2464 53032
rect 2780 53023 2832 53032
rect 2780 52989 2789 53023
rect 2789 52989 2823 53023
rect 2823 52989 2832 53023
rect 2780 52980 2832 52989
rect 26792 52980 26844 53032
rect 23204 52887 23256 52896
rect 23204 52853 23213 52887
rect 23213 52853 23247 52887
rect 23247 52853 23256 52887
rect 23204 52844 23256 52853
rect 23480 52844 23532 52896
rect 26424 52887 26476 52896
rect 26424 52853 26433 52887
rect 26433 52853 26467 52887
rect 26467 52853 26476 52887
rect 26424 52844 26476 52853
rect 27160 52912 27212 52964
rect 27068 52844 27120 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 2412 52683 2464 52692
rect 2412 52649 2421 52683
rect 2421 52649 2455 52683
rect 2455 52649 2464 52683
rect 2412 52640 2464 52649
rect 22100 52572 22152 52624
rect 26884 52615 26936 52624
rect 26884 52581 26893 52615
rect 26893 52581 26927 52615
rect 26927 52581 26936 52615
rect 26884 52572 26936 52581
rect 25044 52504 25096 52556
rect 2320 52479 2372 52488
rect 2320 52445 2329 52479
rect 2329 52445 2363 52479
rect 2363 52445 2372 52479
rect 2320 52436 2372 52445
rect 3148 52479 3200 52488
rect 3148 52445 3157 52479
rect 3157 52445 3191 52479
rect 3191 52445 3200 52479
rect 3148 52436 3200 52445
rect 5172 52436 5224 52488
rect 21916 52436 21968 52488
rect 26976 52436 27028 52488
rect 29000 52436 29052 52488
rect 30196 52436 30248 52488
rect 3884 52343 3936 52352
rect 3884 52309 3893 52343
rect 3893 52309 3927 52343
rect 3927 52309 3936 52343
rect 3884 52300 3936 52309
rect 22468 52368 22520 52420
rect 22652 52300 22704 52352
rect 23756 52300 23808 52352
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 22560 52096 22612 52148
rect 23112 52096 23164 52148
rect 3884 52028 3936 52080
rect 22100 52028 22152 52080
rect 23664 52096 23716 52148
rect 26792 52096 26844 52148
rect 26976 52139 27028 52148
rect 26976 52105 26985 52139
rect 26985 52105 27019 52139
rect 27019 52105 27028 52139
rect 26976 52096 27028 52105
rect 27068 52028 27120 52080
rect 19984 52003 20036 52012
rect 19984 51969 19993 52003
rect 19993 51969 20027 52003
rect 20027 51969 20036 52003
rect 19984 51960 20036 51969
rect 20076 52003 20128 52012
rect 20076 51969 20085 52003
rect 20085 51969 20119 52003
rect 20119 51969 20128 52003
rect 21916 52003 21968 52012
rect 20076 51960 20128 51969
rect 21916 51969 21925 52003
rect 21925 51969 21959 52003
rect 21959 51969 21968 52003
rect 21916 51960 21968 51969
rect 23204 51960 23256 52012
rect 25044 52003 25096 52012
rect 25044 51969 25053 52003
rect 25053 51969 25087 52003
rect 25087 51969 25096 52003
rect 25044 51960 25096 51969
rect 26424 51960 26476 52012
rect 29000 51960 29052 52012
rect 29552 51960 29604 52012
rect 32128 52028 32180 52080
rect 30472 52003 30524 52012
rect 30472 51969 30506 52003
rect 30506 51969 30524 52003
rect 30472 51960 30524 51969
rect 31392 51960 31444 52012
rect 3148 51892 3200 51944
rect 3240 51935 3292 51944
rect 3240 51901 3249 51935
rect 3249 51901 3283 51935
rect 3283 51901 3292 51935
rect 3240 51892 3292 51901
rect 23756 51867 23808 51876
rect 23756 51833 23765 51867
rect 23765 51833 23799 51867
rect 23799 51833 23808 51867
rect 23756 51824 23808 51833
rect 32404 51892 32456 51944
rect 19340 51756 19392 51808
rect 24216 51756 24268 51808
rect 32312 51756 32364 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 22192 51552 22244 51604
rect 22652 51595 22704 51604
rect 22652 51561 22661 51595
rect 22661 51561 22695 51595
rect 22695 51561 22704 51595
rect 22652 51552 22704 51561
rect 23664 51552 23716 51604
rect 27344 51552 27396 51604
rect 30472 51552 30524 51604
rect 19248 51391 19300 51400
rect 19248 51357 19257 51391
rect 19257 51357 19291 51391
rect 19291 51357 19300 51391
rect 19248 51348 19300 51357
rect 19340 51348 19392 51400
rect 22376 51348 22428 51400
rect 22744 51348 22796 51400
rect 23204 51459 23256 51468
rect 23204 51425 23213 51459
rect 23213 51425 23247 51459
rect 23247 51425 23256 51459
rect 23204 51416 23256 51425
rect 26884 51416 26936 51468
rect 23756 51348 23808 51400
rect 25780 51391 25832 51400
rect 25780 51357 25789 51391
rect 25789 51357 25823 51391
rect 25823 51357 25832 51391
rect 25780 51348 25832 51357
rect 29644 51348 29696 51400
rect 29736 51391 29788 51400
rect 29736 51357 29745 51391
rect 29745 51357 29779 51391
rect 29779 51357 29788 51391
rect 29736 51348 29788 51357
rect 23112 51323 23164 51332
rect 23112 51289 23121 51323
rect 23121 51289 23155 51323
rect 23155 51289 23164 51323
rect 23112 51280 23164 51289
rect 25504 51280 25556 51332
rect 31392 51391 31444 51400
rect 31392 51357 31401 51391
rect 31401 51357 31435 51391
rect 31435 51357 31444 51391
rect 31392 51348 31444 51357
rect 32128 51348 32180 51400
rect 32312 51391 32364 51400
rect 32312 51357 32346 51391
rect 32346 51357 32364 51391
rect 32312 51348 32364 51357
rect 32588 51348 32640 51400
rect 36176 51348 36228 51400
rect 57520 51348 57572 51400
rect 57796 51391 57848 51400
rect 57796 51357 57805 51391
rect 57805 51357 57839 51391
rect 57839 51357 57848 51391
rect 57796 51348 57848 51357
rect 32496 51280 32548 51332
rect 33140 51280 33192 51332
rect 20628 51255 20680 51264
rect 20628 51221 20637 51255
rect 20637 51221 20671 51255
rect 20671 51221 20680 51255
rect 20628 51212 20680 51221
rect 24584 51212 24636 51264
rect 28816 51255 28868 51264
rect 28816 51221 28825 51255
rect 28825 51221 28859 51255
rect 28859 51221 28868 51255
rect 28816 51212 28868 51221
rect 33048 51212 33100 51264
rect 33416 51255 33468 51264
rect 33416 51221 33425 51255
rect 33425 51221 33459 51255
rect 33459 51221 33468 51255
rect 33416 51212 33468 51221
rect 33876 51255 33928 51264
rect 33876 51221 33885 51255
rect 33885 51221 33919 51255
rect 33919 51221 33928 51255
rect 33876 51212 33928 51221
rect 57060 51255 57112 51264
rect 57060 51221 57069 51255
rect 57069 51221 57103 51255
rect 57103 51221 57112 51255
rect 57060 51212 57112 51221
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 22468 51008 22520 51060
rect 32588 51008 32640 51060
rect 33140 51008 33192 51060
rect 20260 50940 20312 50992
rect 20628 50940 20680 50992
rect 20076 50872 20128 50924
rect 23204 50940 23256 50992
rect 23480 50915 23532 50924
rect 23480 50881 23489 50915
rect 23489 50881 23523 50915
rect 23523 50881 23532 50915
rect 23480 50872 23532 50881
rect 22744 50804 22796 50856
rect 25504 50872 25556 50924
rect 28264 50872 28316 50924
rect 28908 50940 28960 50992
rect 29460 50940 29512 50992
rect 28816 50915 28868 50924
rect 28816 50881 28850 50915
rect 28850 50881 28868 50915
rect 28816 50872 28868 50881
rect 31392 50915 31444 50924
rect 31392 50881 31401 50915
rect 31401 50881 31435 50915
rect 31435 50881 31444 50915
rect 31392 50872 31444 50881
rect 33876 50940 33928 50992
rect 32680 50872 32732 50924
rect 33324 50872 33376 50924
rect 18696 50668 18748 50720
rect 22376 50668 22428 50720
rect 23480 50736 23532 50788
rect 25596 50804 25648 50856
rect 31668 50804 31720 50856
rect 31944 50804 31996 50856
rect 32128 50847 32180 50856
rect 32128 50813 32137 50847
rect 32137 50813 32171 50847
rect 32171 50813 32180 50847
rect 32128 50804 32180 50813
rect 33508 50804 33560 50856
rect 29828 50736 29880 50788
rect 25780 50668 25832 50720
rect 29736 50668 29788 50720
rect 30840 50668 30892 50720
rect 33968 50711 34020 50720
rect 33968 50677 33977 50711
rect 33977 50677 34011 50711
rect 34011 50677 34020 50711
rect 33968 50668 34020 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 25044 50507 25096 50516
rect 25044 50473 25053 50507
rect 25053 50473 25087 50507
rect 25087 50473 25096 50507
rect 25044 50464 25096 50473
rect 19248 50371 19300 50380
rect 19248 50337 19257 50371
rect 19257 50337 19291 50371
rect 19291 50337 19300 50371
rect 19248 50328 19300 50337
rect 26056 50328 26108 50380
rect 18696 50303 18748 50312
rect 18696 50269 18705 50303
rect 18705 50269 18739 50303
rect 18739 50269 18748 50303
rect 18696 50260 18748 50269
rect 22376 50303 22428 50312
rect 22376 50269 22385 50303
rect 22385 50269 22419 50303
rect 22419 50269 22428 50303
rect 22376 50260 22428 50269
rect 25596 50260 25648 50312
rect 28264 50260 28316 50312
rect 25964 50192 26016 50244
rect 31944 50464 31996 50516
rect 33324 50464 33376 50516
rect 33508 50507 33560 50516
rect 33508 50473 33517 50507
rect 33517 50473 33551 50507
rect 33551 50473 33560 50507
rect 33508 50464 33560 50473
rect 30840 50371 30892 50380
rect 30840 50337 30849 50371
rect 30849 50337 30883 50371
rect 30883 50337 30892 50371
rect 30840 50328 30892 50337
rect 57796 50396 57848 50448
rect 57060 50328 57112 50380
rect 57888 50371 57940 50380
rect 57888 50337 57897 50371
rect 57897 50337 57931 50371
rect 57931 50337 57940 50371
rect 57888 50328 57940 50337
rect 29828 50303 29880 50312
rect 29828 50269 29837 50303
rect 29837 50269 29871 50303
rect 29871 50269 29880 50303
rect 29828 50260 29880 50269
rect 30012 50303 30064 50312
rect 30012 50269 30021 50303
rect 30021 50269 30055 50303
rect 30055 50269 30064 50303
rect 30012 50260 30064 50269
rect 30288 50260 30340 50312
rect 30932 50303 30984 50312
rect 30932 50269 30941 50303
rect 30941 50269 30975 50303
rect 30975 50269 30984 50303
rect 30932 50260 30984 50269
rect 32128 50303 32180 50312
rect 30104 50192 30156 50244
rect 32128 50269 32137 50303
rect 32137 50269 32171 50303
rect 32171 50269 32180 50303
rect 32128 50260 32180 50269
rect 33140 50192 33192 50244
rect 20628 50167 20680 50176
rect 20628 50133 20637 50167
rect 20637 50133 20671 50167
rect 20671 50133 20680 50167
rect 20628 50124 20680 50133
rect 22192 50167 22244 50176
rect 22192 50133 22201 50167
rect 22201 50133 22235 50167
rect 22235 50133 22244 50167
rect 22192 50124 22244 50133
rect 29920 50124 29972 50176
rect 32312 50124 32364 50176
rect 33968 50124 34020 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 19432 49920 19484 49972
rect 19984 49920 20036 49972
rect 20628 49963 20680 49972
rect 20628 49929 20637 49963
rect 20637 49929 20671 49963
rect 20671 49929 20680 49963
rect 20628 49920 20680 49929
rect 29552 49920 29604 49972
rect 30104 49920 30156 49972
rect 30932 49963 30984 49972
rect 30932 49929 30941 49963
rect 30941 49929 30975 49963
rect 30975 49929 30984 49963
rect 30932 49920 30984 49929
rect 32312 49963 32364 49972
rect 32312 49929 32321 49963
rect 32321 49929 32355 49963
rect 32355 49929 32364 49963
rect 32312 49920 32364 49929
rect 32496 49963 32548 49972
rect 32496 49929 32505 49963
rect 32505 49929 32539 49963
rect 32539 49929 32548 49963
rect 32496 49920 32548 49929
rect 32680 49963 32732 49972
rect 32680 49929 32689 49963
rect 32689 49929 32723 49963
rect 32723 49929 32732 49963
rect 32680 49920 32732 49929
rect 33140 49963 33192 49972
rect 33140 49929 33149 49963
rect 33149 49929 33183 49963
rect 33183 49929 33192 49963
rect 33140 49920 33192 49929
rect 20260 49895 20312 49904
rect 20260 49861 20269 49895
rect 20269 49861 20303 49895
rect 20303 49861 20312 49895
rect 20260 49852 20312 49861
rect 24032 49852 24084 49904
rect 27620 49895 27672 49904
rect 27620 49861 27629 49895
rect 27629 49861 27663 49895
rect 27663 49861 27672 49895
rect 27620 49852 27672 49861
rect 20076 49784 20128 49836
rect 20536 49827 20588 49836
rect 20536 49793 20545 49827
rect 20545 49793 20579 49827
rect 20579 49793 20588 49827
rect 20536 49784 20588 49793
rect 3424 49716 3476 49768
rect 9680 49716 9732 49768
rect 20168 49716 20220 49768
rect 20628 49716 20680 49768
rect 22008 49716 22060 49768
rect 23480 49827 23532 49836
rect 23480 49793 23489 49827
rect 23489 49793 23523 49827
rect 23523 49793 23532 49827
rect 23480 49784 23532 49793
rect 24124 49784 24176 49836
rect 24400 49827 24452 49836
rect 24400 49793 24409 49827
rect 24409 49793 24443 49827
rect 24443 49793 24452 49827
rect 24400 49784 24452 49793
rect 28264 49827 28316 49836
rect 28264 49793 28273 49827
rect 28273 49793 28307 49827
rect 28307 49793 28316 49827
rect 28264 49784 28316 49793
rect 31668 49852 31720 49904
rect 33508 49852 33560 49904
rect 29092 49784 29144 49836
rect 29276 49784 29328 49836
rect 33048 49784 33100 49836
rect 37832 49827 37884 49836
rect 37832 49793 37866 49827
rect 37866 49793 37884 49827
rect 37832 49784 37884 49793
rect 39212 49784 39264 49836
rect 39948 49784 40000 49836
rect 40316 49827 40368 49836
rect 40316 49793 40325 49827
rect 40325 49793 40359 49827
rect 40359 49793 40368 49827
rect 40316 49784 40368 49793
rect 23572 49716 23624 49768
rect 23848 49716 23900 49768
rect 24676 49759 24728 49768
rect 24676 49725 24685 49759
rect 24685 49725 24719 49759
rect 24719 49725 24728 49759
rect 24676 49716 24728 49725
rect 25596 49716 25648 49768
rect 25780 49716 25832 49768
rect 30104 49759 30156 49768
rect 30104 49725 30113 49759
rect 30113 49725 30147 49759
rect 30147 49725 30156 49759
rect 30104 49716 30156 49725
rect 37372 49716 37424 49768
rect 39672 49759 39724 49768
rect 39672 49725 39681 49759
rect 39681 49725 39715 49759
rect 39715 49725 39724 49759
rect 39672 49716 39724 49725
rect 41512 49716 41564 49768
rect 23480 49648 23532 49700
rect 22376 49580 22428 49632
rect 38936 49623 38988 49632
rect 38936 49589 38945 49623
rect 38945 49589 38979 49623
rect 38979 49589 38988 49623
rect 38936 49580 38988 49589
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19248 49376 19300 49428
rect 19248 49283 19300 49292
rect 19248 49249 19257 49283
rect 19257 49249 19291 49283
rect 19291 49249 19300 49283
rect 19248 49240 19300 49249
rect 23572 49376 23624 49428
rect 29184 49376 29236 49428
rect 29460 49376 29512 49428
rect 29920 49376 29972 49428
rect 39948 49376 40000 49428
rect 24124 49240 24176 49292
rect 26056 49240 26108 49292
rect 29736 49283 29788 49292
rect 21640 49215 21692 49224
rect 19432 49104 19484 49156
rect 21640 49181 21649 49215
rect 21649 49181 21683 49215
rect 21683 49181 21692 49215
rect 21640 49172 21692 49181
rect 22192 49172 22244 49224
rect 23664 49215 23716 49224
rect 23664 49181 23673 49215
rect 23673 49181 23707 49215
rect 23707 49181 23716 49215
rect 23664 49172 23716 49181
rect 25044 49172 25096 49224
rect 29736 49249 29745 49283
rect 29745 49249 29779 49283
rect 29779 49249 29788 49283
rect 29736 49240 29788 49249
rect 23756 49104 23808 49156
rect 20628 49079 20680 49088
rect 20628 49045 20637 49079
rect 20637 49045 20671 49079
rect 20671 49045 20680 49079
rect 20628 49036 20680 49045
rect 24032 49036 24084 49088
rect 28264 49172 28316 49224
rect 29552 49215 29604 49224
rect 29552 49181 29561 49215
rect 29561 49181 29595 49215
rect 29595 49181 29604 49215
rect 29552 49172 29604 49181
rect 38936 49240 38988 49292
rect 39856 49283 39908 49292
rect 39856 49249 39865 49283
rect 39865 49249 39899 49283
rect 39899 49249 39908 49283
rect 39856 49240 39908 49249
rect 48964 49283 49016 49292
rect 30104 49172 30156 49224
rect 32128 49172 32180 49224
rect 37372 49215 37424 49224
rect 37372 49181 37381 49215
rect 37381 49181 37415 49215
rect 37415 49181 37424 49215
rect 37372 49172 37424 49181
rect 40132 49215 40184 49224
rect 40132 49181 40141 49215
rect 40141 49181 40175 49215
rect 40175 49181 40184 49215
rect 40132 49172 40184 49181
rect 40316 49172 40368 49224
rect 41788 49172 41840 49224
rect 27896 49147 27948 49156
rect 27896 49113 27930 49147
rect 27930 49113 27948 49147
rect 30564 49147 30616 49156
rect 27896 49104 27948 49113
rect 30564 49113 30573 49147
rect 30573 49113 30607 49147
rect 30607 49113 30616 49147
rect 30564 49104 30616 49113
rect 34244 49104 34296 49156
rect 37280 49104 37332 49156
rect 41972 49104 42024 49156
rect 42708 49172 42760 49224
rect 48964 49249 48973 49283
rect 48973 49249 49007 49283
rect 49007 49249 49016 49283
rect 48964 49240 49016 49249
rect 47768 49215 47820 49224
rect 47768 49181 47777 49215
rect 47777 49181 47811 49215
rect 47811 49181 47820 49215
rect 47768 49172 47820 49181
rect 56600 49172 56652 49224
rect 43536 49104 43588 49156
rect 48228 49104 48280 49156
rect 57244 49172 57296 49224
rect 57612 49104 57664 49156
rect 27160 49036 27212 49088
rect 36084 49079 36136 49088
rect 36084 49045 36093 49079
rect 36093 49045 36127 49079
rect 36127 49045 36136 49079
rect 36084 49036 36136 49045
rect 38752 49079 38804 49088
rect 38752 49045 38761 49079
rect 38761 49045 38795 49079
rect 38795 49045 38804 49079
rect 38752 49036 38804 49045
rect 42892 49036 42944 49088
rect 44456 49036 44508 49088
rect 57152 49079 57204 49088
rect 57152 49045 57161 49079
rect 57161 49045 57195 49079
rect 57195 49045 57204 49079
rect 57152 49036 57204 49045
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 23480 48875 23532 48884
rect 23480 48841 23489 48875
rect 23489 48841 23523 48875
rect 23523 48841 23532 48875
rect 23480 48832 23532 48841
rect 24308 48832 24360 48884
rect 19156 48764 19208 48816
rect 20168 48807 20220 48816
rect 20168 48773 20177 48807
rect 20177 48773 20211 48807
rect 20211 48773 20220 48807
rect 20168 48764 20220 48773
rect 20260 48764 20312 48816
rect 21640 48764 21692 48816
rect 27896 48832 27948 48884
rect 34244 48875 34296 48884
rect 34244 48841 34253 48875
rect 34253 48841 34287 48875
rect 34287 48841 34296 48875
rect 34244 48832 34296 48841
rect 36084 48832 36136 48884
rect 47768 48832 47820 48884
rect 48228 48875 48280 48884
rect 48228 48841 48237 48875
rect 48237 48841 48271 48875
rect 48271 48841 48280 48875
rect 48228 48832 48280 48841
rect 22376 48739 22428 48748
rect 22376 48705 22410 48739
rect 22410 48705 22428 48739
rect 22376 48696 22428 48705
rect 24032 48739 24084 48748
rect 24032 48705 24041 48739
rect 24041 48705 24075 48739
rect 24075 48705 24084 48739
rect 24032 48696 24084 48705
rect 24308 48739 24360 48748
rect 24308 48705 24317 48739
rect 24317 48705 24351 48739
rect 24351 48705 24360 48739
rect 24308 48696 24360 48705
rect 25044 48739 25096 48748
rect 25044 48705 25053 48739
rect 25053 48705 25087 48739
rect 25087 48705 25096 48739
rect 25044 48696 25096 48705
rect 27160 48739 27212 48748
rect 27160 48705 27169 48739
rect 27169 48705 27203 48739
rect 27203 48705 27212 48739
rect 27160 48696 27212 48705
rect 28080 48696 28132 48748
rect 29368 48764 29420 48816
rect 29644 48807 29696 48816
rect 29644 48773 29653 48807
rect 29653 48773 29687 48807
rect 29687 48773 29696 48807
rect 29644 48764 29696 48773
rect 31944 48764 31996 48816
rect 41788 48807 41840 48816
rect 41788 48773 41797 48807
rect 41797 48773 41831 48807
rect 41831 48773 41840 48807
rect 41788 48764 41840 48773
rect 29460 48745 29512 48754
rect 29460 48711 29469 48745
rect 29469 48711 29503 48745
rect 29503 48711 29512 48745
rect 33692 48739 33744 48748
rect 29460 48702 29512 48711
rect 33692 48705 33701 48739
rect 33701 48705 33735 48739
rect 33735 48705 33744 48739
rect 33692 48696 33744 48705
rect 37372 48739 37424 48748
rect 8484 48671 8536 48680
rect 8484 48637 8493 48671
rect 8493 48637 8527 48671
rect 8527 48637 8536 48671
rect 8484 48628 8536 48637
rect 9680 48671 9732 48680
rect 9680 48637 9689 48671
rect 9689 48637 9723 48671
rect 9723 48637 9732 48671
rect 9680 48628 9732 48637
rect 19708 48628 19760 48680
rect 20628 48628 20680 48680
rect 24400 48628 24452 48680
rect 19984 48492 20036 48544
rect 21364 48492 21416 48544
rect 24124 48535 24176 48544
rect 24124 48501 24133 48535
rect 24133 48501 24167 48535
rect 24167 48501 24176 48535
rect 24124 48492 24176 48501
rect 24400 48492 24452 48544
rect 29000 48560 29052 48612
rect 29184 48560 29236 48612
rect 32588 48628 32640 48680
rect 37372 48705 37381 48739
rect 37381 48705 37415 48739
rect 37415 48705 37424 48739
rect 37372 48696 37424 48705
rect 38200 48696 38252 48748
rect 38752 48696 38804 48748
rect 39948 48696 40000 48748
rect 41880 48739 41932 48748
rect 39212 48671 39264 48680
rect 39212 48637 39221 48671
rect 39221 48637 39255 48671
rect 39255 48637 39264 48671
rect 39212 48628 39264 48637
rect 29552 48560 29604 48612
rect 40132 48628 40184 48680
rect 40592 48628 40644 48680
rect 41144 48628 41196 48680
rect 41880 48705 41889 48739
rect 41889 48705 41923 48739
rect 41923 48705 41932 48739
rect 41880 48696 41932 48705
rect 44916 48739 44968 48748
rect 42524 48628 42576 48680
rect 42708 48628 42760 48680
rect 44916 48705 44925 48739
rect 44925 48705 44959 48739
rect 44959 48705 44968 48739
rect 44916 48696 44968 48705
rect 45008 48739 45060 48748
rect 45008 48705 45017 48739
rect 45017 48705 45051 48739
rect 45051 48705 45060 48739
rect 45008 48696 45060 48705
rect 45192 48696 45244 48748
rect 48136 48739 48188 48748
rect 48136 48705 48145 48739
rect 48145 48705 48179 48739
rect 48179 48705 48188 48739
rect 48136 48696 48188 48705
rect 56876 48696 56928 48748
rect 41880 48560 41932 48612
rect 46020 48628 46072 48680
rect 40684 48492 40736 48544
rect 43996 48535 44048 48544
rect 43996 48501 44005 48535
rect 44005 48501 44039 48535
rect 44039 48501 44048 48535
rect 43996 48492 44048 48501
rect 45284 48535 45336 48544
rect 45284 48501 45293 48535
rect 45293 48501 45327 48535
rect 45327 48501 45336 48535
rect 45284 48492 45336 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 23756 48288 23808 48340
rect 37280 48331 37332 48340
rect 37280 48297 37289 48331
rect 37289 48297 37323 48331
rect 37323 48297 37332 48331
rect 37280 48288 37332 48297
rect 38200 48288 38252 48340
rect 26976 48220 27028 48272
rect 30196 48220 30248 48272
rect 25596 48195 25648 48204
rect 25596 48161 25605 48195
rect 25605 48161 25639 48195
rect 25639 48161 25648 48195
rect 25596 48152 25648 48161
rect 28080 48195 28132 48204
rect 28080 48161 28089 48195
rect 28089 48161 28123 48195
rect 28123 48161 28132 48195
rect 28080 48152 28132 48161
rect 19708 48127 19760 48136
rect 19708 48093 19717 48127
rect 19717 48093 19751 48127
rect 19751 48093 19760 48127
rect 19708 48084 19760 48093
rect 19984 48084 20036 48136
rect 23848 48127 23900 48136
rect 23848 48093 23857 48127
rect 23857 48093 23891 48127
rect 23891 48093 23900 48127
rect 23848 48084 23900 48093
rect 24400 48127 24452 48136
rect 24400 48093 24409 48127
rect 24409 48093 24443 48127
rect 24443 48093 24452 48127
rect 24400 48084 24452 48093
rect 24584 48127 24636 48136
rect 24584 48093 24593 48127
rect 24593 48093 24627 48127
rect 24627 48093 24636 48127
rect 24584 48084 24636 48093
rect 26148 48084 26200 48136
rect 27620 48084 27672 48136
rect 29276 48084 29328 48136
rect 31024 48084 31076 48136
rect 34152 48084 34204 48136
rect 36544 48084 36596 48136
rect 39764 48220 39816 48272
rect 37188 48084 37240 48136
rect 38108 48127 38160 48136
rect 38108 48093 38117 48127
rect 38117 48093 38151 48127
rect 38151 48093 38160 48127
rect 38108 48084 38160 48093
rect 39948 48127 40000 48136
rect 39948 48093 39957 48127
rect 39957 48093 39991 48127
rect 39991 48093 40000 48127
rect 39948 48084 40000 48093
rect 40592 48127 40644 48136
rect 40592 48093 40601 48127
rect 40601 48093 40635 48127
rect 40635 48093 40644 48127
rect 40592 48084 40644 48093
rect 41880 48288 41932 48340
rect 46020 48331 46072 48340
rect 46020 48297 46029 48331
rect 46029 48297 46063 48331
rect 46063 48297 46072 48331
rect 46020 48288 46072 48297
rect 40960 48220 41012 48272
rect 45284 48220 45336 48272
rect 41052 48195 41104 48204
rect 41052 48161 41061 48195
rect 41061 48161 41095 48195
rect 41095 48161 41104 48195
rect 41052 48152 41104 48161
rect 41788 48152 41840 48204
rect 41144 48127 41196 48136
rect 19156 48016 19208 48068
rect 30472 48016 30524 48068
rect 31944 48059 31996 48068
rect 31944 48025 31953 48059
rect 31953 48025 31987 48059
rect 31987 48025 31996 48059
rect 31944 48016 31996 48025
rect 33048 48059 33100 48068
rect 33048 48025 33082 48059
rect 33082 48025 33100 48059
rect 20812 47948 20864 48000
rect 24768 47991 24820 48000
rect 24768 47957 24777 47991
rect 24777 47957 24811 47991
rect 24811 47957 24820 47991
rect 24768 47948 24820 47957
rect 31760 47948 31812 48000
rect 33048 48016 33100 48025
rect 33324 47948 33376 48000
rect 33692 47948 33744 48000
rect 37372 47948 37424 48000
rect 39672 48016 39724 48068
rect 41144 48093 41153 48127
rect 41153 48093 41187 48127
rect 41187 48093 41196 48127
rect 41144 48084 41196 48093
rect 40868 48016 40920 48068
rect 41972 48084 42024 48136
rect 44088 48152 44140 48204
rect 44272 48152 44324 48204
rect 48136 48220 48188 48272
rect 43996 48084 44048 48136
rect 45192 48127 45244 48136
rect 45192 48093 45201 48127
rect 45201 48093 45235 48127
rect 45235 48093 45244 48127
rect 45192 48084 45244 48093
rect 42892 48016 42944 48068
rect 45376 48084 45428 48136
rect 46572 48152 46624 48204
rect 57244 48220 57296 48272
rect 57152 48152 57204 48204
rect 57888 48195 57940 48204
rect 57888 48161 57897 48195
rect 57897 48161 57931 48195
rect 57931 48161 57940 48195
rect 57888 48152 57940 48161
rect 46296 48127 46348 48136
rect 45836 48016 45888 48068
rect 46296 48093 46305 48127
rect 46305 48093 46339 48127
rect 46339 48093 46348 48127
rect 46296 48084 46348 48093
rect 46388 48016 46440 48068
rect 46940 48016 46992 48068
rect 47400 48084 47452 48136
rect 47676 48016 47728 48068
rect 43628 47948 43680 48000
rect 45468 47948 45520 48000
rect 46204 47991 46256 48000
rect 46204 47957 46213 47991
rect 46213 47957 46247 47991
rect 46247 47957 46256 47991
rect 46204 47948 46256 47957
rect 47768 47948 47820 48000
rect 48780 47948 48832 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 24676 47744 24728 47796
rect 33048 47787 33100 47796
rect 33048 47753 33057 47787
rect 33057 47753 33091 47787
rect 33091 47753 33100 47787
rect 33048 47744 33100 47753
rect 33876 47744 33928 47796
rect 37832 47787 37884 47796
rect 24768 47676 24820 47728
rect 29552 47676 29604 47728
rect 30564 47676 30616 47728
rect 37556 47719 37608 47728
rect 8944 47608 8996 47660
rect 20812 47651 20864 47660
rect 18788 47583 18840 47592
rect 18788 47549 18797 47583
rect 18797 47549 18831 47583
rect 18831 47549 18840 47583
rect 18788 47540 18840 47549
rect 20812 47617 20821 47651
rect 20821 47617 20855 47651
rect 20855 47617 20864 47651
rect 20812 47608 20864 47617
rect 24216 47651 24268 47660
rect 24216 47617 24225 47651
rect 24225 47617 24259 47651
rect 24259 47617 24268 47651
rect 24216 47608 24268 47617
rect 26056 47608 26108 47660
rect 26148 47608 26200 47660
rect 27620 47651 27672 47660
rect 27620 47617 27629 47651
rect 27629 47617 27663 47651
rect 27663 47617 27672 47651
rect 27620 47608 27672 47617
rect 28264 47651 28316 47660
rect 28264 47617 28273 47651
rect 28273 47617 28307 47651
rect 28307 47617 28316 47651
rect 28264 47608 28316 47617
rect 30380 47651 30432 47660
rect 30380 47617 30389 47651
rect 30389 47617 30423 47651
rect 30423 47617 30432 47651
rect 30380 47608 30432 47617
rect 24676 47583 24728 47592
rect 24676 47549 24685 47583
rect 24685 47549 24719 47583
rect 24719 47549 24728 47583
rect 24676 47540 24728 47549
rect 28908 47583 28960 47592
rect 28908 47549 28917 47583
rect 28917 47549 28951 47583
rect 28951 47549 28960 47583
rect 28908 47540 28960 47549
rect 30472 47540 30524 47592
rect 31944 47608 31996 47660
rect 32404 47608 32456 47660
rect 32588 47651 32640 47660
rect 32588 47617 32597 47651
rect 32597 47617 32631 47651
rect 32631 47617 32640 47651
rect 33324 47651 33376 47660
rect 32588 47608 32640 47617
rect 33324 47617 33333 47651
rect 33333 47617 33367 47651
rect 33367 47617 33376 47651
rect 33324 47608 33376 47617
rect 33508 47651 33560 47660
rect 33508 47617 33517 47651
rect 33517 47617 33551 47651
rect 33551 47617 33560 47651
rect 33692 47651 33744 47660
rect 33508 47608 33560 47617
rect 33692 47617 33701 47651
rect 33701 47617 33735 47651
rect 33735 47617 33744 47651
rect 33692 47608 33744 47617
rect 34152 47651 34204 47660
rect 34152 47617 34161 47651
rect 34161 47617 34195 47651
rect 34195 47617 34204 47651
rect 34152 47608 34204 47617
rect 37556 47685 37565 47719
rect 37565 47685 37599 47719
rect 37599 47685 37608 47719
rect 37556 47676 37608 47685
rect 37280 47651 37332 47660
rect 37280 47617 37289 47651
rect 37289 47617 37323 47651
rect 37323 47617 37332 47651
rect 37280 47608 37332 47617
rect 37372 47608 37424 47660
rect 37832 47753 37841 47787
rect 37841 47753 37875 47787
rect 37875 47753 37884 47787
rect 37832 47744 37884 47753
rect 40592 47719 40644 47728
rect 40592 47685 40601 47719
rect 40601 47685 40635 47719
rect 40635 47685 40644 47719
rect 40592 47676 40644 47685
rect 44916 47744 44968 47796
rect 45192 47744 45244 47796
rect 46112 47744 46164 47796
rect 46940 47744 46992 47796
rect 44088 47676 44140 47728
rect 38108 47608 38160 47660
rect 39212 47608 39264 47660
rect 41144 47608 41196 47660
rect 41420 47608 41472 47660
rect 44180 47651 44232 47660
rect 44180 47617 44189 47651
rect 44189 47617 44223 47651
rect 44223 47617 44232 47651
rect 44180 47608 44232 47617
rect 19524 47404 19576 47456
rect 20168 47447 20220 47456
rect 20168 47413 20177 47447
rect 20177 47413 20211 47447
rect 20211 47413 20220 47447
rect 20168 47404 20220 47413
rect 24492 47404 24544 47456
rect 25964 47447 26016 47456
rect 25964 47413 25973 47447
rect 25973 47413 26007 47447
rect 26007 47413 26016 47447
rect 25964 47404 26016 47413
rect 27620 47404 27672 47456
rect 31852 47404 31904 47456
rect 44272 47540 44324 47592
rect 44916 47608 44968 47660
rect 45376 47651 45428 47660
rect 45376 47617 45385 47651
rect 45385 47617 45419 47651
rect 45419 47617 45428 47651
rect 45376 47608 45428 47617
rect 45468 47651 45520 47660
rect 45468 47617 45477 47651
rect 45477 47617 45511 47651
rect 45511 47617 45520 47651
rect 45652 47651 45704 47660
rect 45468 47608 45520 47617
rect 45652 47617 45661 47651
rect 45661 47617 45695 47651
rect 45695 47617 45704 47651
rect 45652 47608 45704 47617
rect 46204 47608 46256 47660
rect 46572 47651 46624 47660
rect 46572 47617 46581 47651
rect 46581 47617 46615 47651
rect 46615 47617 46624 47651
rect 46572 47608 46624 47617
rect 47860 47651 47912 47660
rect 47860 47617 47869 47651
rect 47869 47617 47903 47651
rect 47903 47617 47912 47651
rect 47860 47608 47912 47617
rect 48228 47651 48280 47660
rect 46112 47583 46164 47592
rect 46112 47549 46121 47583
rect 46121 47549 46155 47583
rect 46155 47549 46164 47583
rect 46112 47540 46164 47549
rect 47032 47540 47084 47592
rect 47768 47540 47820 47592
rect 48228 47617 48237 47651
rect 48237 47617 48271 47651
rect 48271 47617 48280 47651
rect 48228 47608 48280 47617
rect 48412 47608 48464 47660
rect 48780 47583 48832 47592
rect 48780 47549 48789 47583
rect 48789 47549 48823 47583
rect 48823 47549 48832 47583
rect 48780 47540 48832 47549
rect 35440 47472 35492 47524
rect 39856 47515 39908 47524
rect 39856 47481 39865 47515
rect 39865 47481 39899 47515
rect 39899 47481 39908 47515
rect 39856 47472 39908 47481
rect 44180 47472 44232 47524
rect 46296 47515 46348 47524
rect 46296 47481 46305 47515
rect 46305 47481 46339 47515
rect 46339 47481 46348 47515
rect 46296 47472 46348 47481
rect 35532 47447 35584 47456
rect 35532 47413 35541 47447
rect 35541 47413 35575 47447
rect 35575 47413 35584 47447
rect 35532 47404 35584 47413
rect 37556 47404 37608 47456
rect 40868 47404 40920 47456
rect 41696 47447 41748 47456
rect 41696 47413 41705 47447
rect 41705 47413 41739 47447
rect 41739 47413 41748 47447
rect 41696 47404 41748 47413
rect 45928 47404 45980 47456
rect 46112 47404 46164 47456
rect 46572 47404 46624 47456
rect 48780 47404 48832 47456
rect 48872 47404 48924 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 2964 47200 3016 47252
rect 19524 47107 19576 47116
rect 19524 47073 19533 47107
rect 19533 47073 19567 47107
rect 19567 47073 19576 47107
rect 19524 47064 19576 47073
rect 20076 47064 20128 47116
rect 19340 46996 19392 47048
rect 19984 46996 20036 47048
rect 20352 47039 20404 47048
rect 19432 46928 19484 46980
rect 20352 47005 20361 47039
rect 20361 47005 20395 47039
rect 20395 47005 20404 47039
rect 20352 46996 20404 47005
rect 21364 47039 21416 47048
rect 21364 47005 21373 47039
rect 21373 47005 21407 47039
rect 21407 47005 21416 47039
rect 21364 46996 21416 47005
rect 24032 46996 24084 47048
rect 20628 46928 20680 46980
rect 22284 46928 22336 46980
rect 27620 47064 27672 47116
rect 40960 47200 41012 47252
rect 41328 47200 41380 47252
rect 30012 47175 30064 47184
rect 30012 47141 30021 47175
rect 30021 47141 30055 47175
rect 30055 47141 30064 47175
rect 30012 47132 30064 47141
rect 30288 47132 30340 47184
rect 31024 47175 31076 47184
rect 31024 47141 31033 47175
rect 31033 47141 31067 47175
rect 31067 47141 31076 47175
rect 31024 47132 31076 47141
rect 35072 47132 35124 47184
rect 37280 47132 37332 47184
rect 37648 47132 37700 47184
rect 39764 47132 39816 47184
rect 45376 47200 45428 47252
rect 47952 47243 48004 47252
rect 47952 47209 47961 47243
rect 47961 47209 47995 47243
rect 47995 47209 48004 47243
rect 47952 47200 48004 47209
rect 48228 47243 48280 47252
rect 48228 47209 48237 47243
rect 48237 47209 48271 47243
rect 48271 47209 48280 47243
rect 48228 47200 48280 47209
rect 30104 47107 30156 47116
rect 30104 47073 30113 47107
rect 30113 47073 30147 47107
rect 30147 47073 30156 47107
rect 30104 47064 30156 47073
rect 30656 47064 30708 47116
rect 31852 47107 31904 47116
rect 31852 47073 31861 47107
rect 31861 47073 31895 47107
rect 31895 47073 31904 47107
rect 31852 47064 31904 47073
rect 33508 47107 33560 47116
rect 33508 47073 33517 47107
rect 33517 47073 33551 47107
rect 33551 47073 33560 47107
rect 33508 47064 33560 47073
rect 35440 47064 35492 47116
rect 41328 47064 41380 47116
rect 24400 47039 24452 47048
rect 24400 47005 24409 47039
rect 24409 47005 24443 47039
rect 24443 47005 24452 47039
rect 24400 46996 24452 47005
rect 24492 46996 24544 47048
rect 26148 46996 26200 47048
rect 27160 47039 27212 47048
rect 27160 47005 27169 47039
rect 27169 47005 27203 47039
rect 27203 47005 27212 47039
rect 27160 46996 27212 47005
rect 30564 46996 30616 47048
rect 35072 47039 35124 47048
rect 35072 47005 35081 47039
rect 35081 47005 35115 47039
rect 35115 47005 35124 47039
rect 35072 46996 35124 47005
rect 27620 46928 27672 46980
rect 31392 46928 31444 46980
rect 33600 46928 33652 46980
rect 22652 46903 22704 46912
rect 22652 46869 22661 46903
rect 22661 46869 22695 46903
rect 22695 46869 22704 46903
rect 22652 46860 22704 46869
rect 25780 46903 25832 46912
rect 25780 46869 25789 46903
rect 25789 46869 25823 46903
rect 25823 46869 25832 46903
rect 25780 46860 25832 46869
rect 26976 46860 27028 46912
rect 34704 46860 34756 46912
rect 35900 46996 35952 47048
rect 35532 46928 35584 46980
rect 39672 46996 39724 47048
rect 39764 46996 39816 47048
rect 37924 46928 37976 46980
rect 40316 47039 40368 47048
rect 40316 47005 40325 47039
rect 40325 47005 40359 47039
rect 40359 47005 40368 47039
rect 41420 47039 41472 47048
rect 40316 46996 40368 47005
rect 41420 47005 41429 47039
rect 41429 47005 41463 47039
rect 41463 47005 41472 47039
rect 56232 47132 56284 47184
rect 44916 47064 44968 47116
rect 41420 46996 41472 47005
rect 42892 46996 42944 47048
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 45376 46996 45428 47048
rect 41972 46928 42024 46980
rect 40316 46903 40368 46912
rect 40316 46869 40325 46903
rect 40325 46869 40359 46903
rect 40359 46869 40368 46903
rect 40316 46860 40368 46869
rect 41512 46860 41564 46912
rect 42432 46928 42484 46980
rect 42800 46928 42852 46980
rect 44180 46928 44232 46980
rect 45928 46996 45980 47048
rect 46940 47039 46992 47048
rect 46940 47005 46949 47039
rect 46949 47005 46983 47039
rect 46983 47005 46992 47039
rect 46940 46996 46992 47005
rect 47124 47039 47176 47048
rect 47124 47005 47133 47039
rect 47133 47005 47167 47039
rect 47167 47005 47176 47039
rect 47124 46996 47176 47005
rect 47216 47039 47268 47048
rect 47216 47005 47225 47039
rect 47225 47005 47259 47039
rect 47259 47005 47268 47039
rect 47676 47039 47728 47048
rect 47216 46996 47268 47005
rect 47676 47005 47685 47039
rect 47685 47005 47719 47039
rect 47719 47005 47728 47039
rect 47676 46996 47728 47005
rect 47860 46996 47912 47048
rect 48872 47039 48924 47048
rect 48872 47005 48881 47039
rect 48881 47005 48915 47039
rect 48915 47005 48924 47039
rect 48872 46996 48924 47005
rect 58072 47064 58124 47116
rect 49884 46996 49936 47048
rect 49976 46996 50028 47048
rect 45744 46928 45796 46980
rect 47768 46928 47820 46980
rect 43168 46903 43220 46912
rect 43168 46869 43177 46903
rect 43177 46869 43211 46903
rect 43211 46869 43220 46903
rect 43168 46860 43220 46869
rect 44732 46860 44784 46912
rect 46388 46860 46440 46912
rect 48320 46928 48372 46980
rect 49792 46928 49844 46980
rect 56968 46928 57020 46980
rect 58164 46971 58216 46980
rect 58164 46937 58173 46971
rect 58173 46937 58207 46971
rect 58207 46937 58216 46971
rect 58164 46928 58216 46937
rect 48688 46903 48740 46912
rect 48688 46869 48697 46903
rect 48697 46869 48731 46903
rect 48731 46869 48740 46903
rect 48688 46860 48740 46869
rect 49608 46860 49660 46912
rect 49976 46860 50028 46912
rect 50068 46860 50120 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 24032 46699 24084 46708
rect 19984 46588 20036 46640
rect 22284 46631 22336 46640
rect 22284 46597 22319 46631
rect 22319 46597 22336 46631
rect 22284 46588 22336 46597
rect 18788 46520 18840 46572
rect 22008 46563 22060 46572
rect 22008 46529 22017 46563
rect 22017 46529 22051 46563
rect 22051 46529 22060 46563
rect 22008 46520 22060 46529
rect 22100 46563 22152 46572
rect 22100 46529 22109 46563
rect 22109 46529 22143 46563
rect 22143 46529 22152 46563
rect 22100 46520 22152 46529
rect 22652 46520 22704 46572
rect 24032 46665 24041 46699
rect 24041 46665 24075 46699
rect 24075 46665 24084 46699
rect 24032 46656 24084 46665
rect 24860 46656 24912 46708
rect 26148 46656 26200 46708
rect 27620 46699 27672 46708
rect 27620 46665 27629 46699
rect 27629 46665 27663 46699
rect 27663 46665 27672 46699
rect 27620 46656 27672 46665
rect 30012 46656 30064 46708
rect 31392 46699 31444 46708
rect 31392 46665 31401 46699
rect 31401 46665 31435 46699
rect 31435 46665 31444 46699
rect 31392 46656 31444 46665
rect 25964 46588 26016 46640
rect 27712 46588 27764 46640
rect 24860 46520 24912 46572
rect 28264 46563 28316 46572
rect 28264 46529 28273 46563
rect 28273 46529 28307 46563
rect 28307 46529 28316 46563
rect 28264 46520 28316 46529
rect 31024 46588 31076 46640
rect 30288 46563 30340 46572
rect 30288 46529 30322 46563
rect 30322 46529 30340 46563
rect 30288 46520 30340 46529
rect 23664 46495 23716 46504
rect 23664 46461 23673 46495
rect 23673 46461 23707 46495
rect 23707 46461 23716 46495
rect 23664 46452 23716 46461
rect 25136 46452 25188 46504
rect 25780 46452 25832 46504
rect 25964 46452 26016 46504
rect 27160 46452 27212 46504
rect 29920 46452 29972 46504
rect 26424 46427 26476 46436
rect 26424 46393 26433 46427
rect 26433 46393 26467 46427
rect 26467 46393 26476 46427
rect 26424 46384 26476 46393
rect 20444 46359 20496 46368
rect 20444 46325 20453 46359
rect 20453 46325 20487 46359
rect 20487 46325 20496 46359
rect 20444 46316 20496 46325
rect 21824 46359 21876 46368
rect 21824 46325 21833 46359
rect 21833 46325 21867 46359
rect 21867 46325 21876 46359
rect 21824 46316 21876 46325
rect 23112 46359 23164 46368
rect 23112 46325 23121 46359
rect 23121 46325 23155 46359
rect 23155 46325 23164 46359
rect 23112 46316 23164 46325
rect 24952 46359 25004 46368
rect 24952 46325 24961 46359
rect 24961 46325 24995 46359
rect 24995 46325 25004 46359
rect 24952 46316 25004 46325
rect 29920 46316 29972 46368
rect 36176 46656 36228 46708
rect 33416 46588 33468 46640
rect 35348 46588 35400 46640
rect 39304 46656 39356 46708
rect 41052 46656 41104 46708
rect 43352 46656 43404 46708
rect 45100 46699 45152 46708
rect 45100 46665 45109 46699
rect 45109 46665 45143 46699
rect 45143 46665 45152 46699
rect 45100 46656 45152 46665
rect 50068 46656 50120 46708
rect 56968 46699 57020 46708
rect 56968 46665 56977 46699
rect 56977 46665 57011 46699
rect 57011 46665 57020 46699
rect 56968 46656 57020 46665
rect 32404 46563 32456 46572
rect 32404 46529 32413 46563
rect 32413 46529 32447 46563
rect 32447 46529 32456 46563
rect 32404 46520 32456 46529
rect 32128 46359 32180 46368
rect 32128 46325 32137 46359
rect 32137 46325 32171 46359
rect 32171 46325 32180 46359
rect 32128 46316 32180 46325
rect 33600 46520 33652 46572
rect 34704 46520 34756 46572
rect 37280 46520 37332 46572
rect 37924 46563 37976 46572
rect 37924 46529 37933 46563
rect 37933 46529 37967 46563
rect 37967 46529 37976 46563
rect 37924 46520 37976 46529
rect 39212 46563 39264 46572
rect 32588 46384 32640 46436
rect 35900 46452 35952 46504
rect 39212 46529 39221 46563
rect 39221 46529 39255 46563
rect 39255 46529 39264 46563
rect 39212 46520 39264 46529
rect 39764 46520 39816 46572
rect 40132 46563 40184 46572
rect 40132 46529 40141 46563
rect 40141 46529 40175 46563
rect 40175 46529 40184 46563
rect 40132 46520 40184 46529
rect 40316 46563 40368 46572
rect 40316 46529 40325 46563
rect 40325 46529 40359 46563
rect 40359 46529 40368 46563
rect 40316 46520 40368 46529
rect 40868 46520 40920 46572
rect 42248 46520 42300 46572
rect 42892 46588 42944 46640
rect 44732 46631 44784 46640
rect 42800 46520 42852 46572
rect 44732 46597 44741 46631
rect 44741 46597 44775 46631
rect 44775 46597 44784 46631
rect 44732 46588 44784 46597
rect 48688 46588 48740 46640
rect 43628 46563 43680 46572
rect 43628 46529 43637 46563
rect 43637 46529 43671 46563
rect 43671 46529 43680 46563
rect 43904 46563 43956 46572
rect 43628 46520 43680 46529
rect 43904 46529 43913 46563
rect 43913 46529 43947 46563
rect 43947 46529 43956 46563
rect 43904 46520 43956 46529
rect 45192 46520 45244 46572
rect 45560 46563 45612 46572
rect 45560 46529 45569 46563
rect 45569 46529 45603 46563
rect 45603 46529 45612 46563
rect 45560 46520 45612 46529
rect 45744 46563 45796 46572
rect 45744 46529 45753 46563
rect 45753 46529 45787 46563
rect 45787 46529 45796 46563
rect 45744 46520 45796 46529
rect 46848 46563 46900 46572
rect 46848 46529 46857 46563
rect 46857 46529 46891 46563
rect 46891 46529 46900 46563
rect 46848 46520 46900 46529
rect 49792 46520 49844 46572
rect 50068 46563 50120 46572
rect 50068 46529 50077 46563
rect 50077 46529 50111 46563
rect 50111 46529 50120 46563
rect 50068 46520 50120 46529
rect 50712 46563 50764 46572
rect 50712 46529 50721 46563
rect 50721 46529 50755 46563
rect 50755 46529 50764 46563
rect 50712 46520 50764 46529
rect 58072 46563 58124 46572
rect 41052 46452 41104 46504
rect 44180 46452 44232 46504
rect 45284 46452 45336 46504
rect 46204 46452 46256 46504
rect 47676 46452 47728 46504
rect 47768 46452 47820 46504
rect 51264 46452 51316 46504
rect 38844 46384 38896 46436
rect 58072 46529 58081 46563
rect 58081 46529 58115 46563
rect 58115 46529 58124 46563
rect 58072 46520 58124 46529
rect 36728 46316 36780 46368
rect 38476 46316 38528 46368
rect 39304 46316 39356 46368
rect 42708 46316 42760 46368
rect 48412 46316 48464 46368
rect 49884 46359 49936 46368
rect 49884 46325 49893 46359
rect 49893 46325 49927 46359
rect 49927 46325 49936 46359
rect 49884 46316 49936 46325
rect 50988 46316 51040 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 20536 46112 20588 46164
rect 26056 46112 26108 46164
rect 29000 46155 29052 46164
rect 20260 46044 20312 46096
rect 23664 46044 23716 46096
rect 24216 46044 24268 46096
rect 29000 46121 29009 46155
rect 29009 46121 29043 46155
rect 29043 46121 29052 46155
rect 29000 46112 29052 46121
rect 33416 46112 33468 46164
rect 33692 46112 33744 46164
rect 18788 45976 18840 46028
rect 19156 45908 19208 45960
rect 24400 46019 24452 46028
rect 19340 45840 19392 45892
rect 22376 45908 22428 45960
rect 23112 45908 23164 45960
rect 24400 45985 24409 46019
rect 24409 45985 24443 46019
rect 24443 45985 24452 46019
rect 24400 45976 24452 45985
rect 29736 45976 29788 46028
rect 30380 45976 30432 46028
rect 31024 46019 31076 46028
rect 31024 45985 31033 46019
rect 31033 45985 31067 46019
rect 31067 45985 31076 46019
rect 31024 45976 31076 45985
rect 24952 45908 25004 45960
rect 27620 45951 27672 45960
rect 27620 45917 27629 45951
rect 27629 45917 27663 45951
rect 27663 45917 27672 45951
rect 27620 45908 27672 45917
rect 28264 45908 28316 45960
rect 32128 45908 32180 45960
rect 35808 46044 35860 46096
rect 33784 45951 33836 45960
rect 21824 45840 21876 45892
rect 24676 45883 24728 45892
rect 24676 45849 24710 45883
rect 24710 45849 24728 45883
rect 24676 45840 24728 45849
rect 26976 45883 27028 45892
rect 26976 45849 26985 45883
rect 26985 45849 27019 45883
rect 27019 45849 27028 45883
rect 26976 45840 27028 45849
rect 27712 45840 27764 45892
rect 25596 45772 25648 45824
rect 32588 45772 32640 45824
rect 33140 45815 33192 45824
rect 33140 45781 33149 45815
rect 33149 45781 33183 45815
rect 33183 45781 33192 45815
rect 33140 45772 33192 45781
rect 33784 45917 33793 45951
rect 33793 45917 33827 45951
rect 33827 45917 33836 45951
rect 33784 45908 33836 45917
rect 34888 45951 34940 45960
rect 33692 45840 33744 45892
rect 34888 45917 34897 45951
rect 34897 45917 34931 45951
rect 34931 45917 34940 45951
rect 34888 45908 34940 45917
rect 35992 45951 36044 45960
rect 35992 45917 36001 45951
rect 36001 45917 36035 45951
rect 36035 45917 36044 45951
rect 35992 45908 36044 45917
rect 37004 45908 37056 45960
rect 37832 45908 37884 45960
rect 38384 46112 38436 46164
rect 42708 46112 42760 46164
rect 45008 46112 45060 46164
rect 45744 46112 45796 46164
rect 47768 46155 47820 46164
rect 47768 46121 47777 46155
rect 47777 46121 47811 46155
rect 47811 46121 47820 46155
rect 47768 46112 47820 46121
rect 47952 46155 48004 46164
rect 47952 46121 47961 46155
rect 47961 46121 47995 46155
rect 47995 46121 48004 46155
rect 47952 46112 48004 46121
rect 38108 45951 38160 45960
rect 38108 45917 38117 45951
rect 38117 45917 38151 45951
rect 38151 45917 38160 45951
rect 38108 45908 38160 45917
rect 38476 45908 38528 45960
rect 39120 45976 39172 46028
rect 38936 45951 38988 45960
rect 38936 45917 38945 45951
rect 38945 45917 38979 45951
rect 38979 45917 38988 45951
rect 38936 45908 38988 45917
rect 41236 46044 41288 46096
rect 43168 46044 43220 46096
rect 45560 46044 45612 46096
rect 49884 46044 49936 46096
rect 37188 45840 37240 45892
rect 38752 45883 38804 45892
rect 38752 45849 38761 45883
rect 38761 45849 38795 45883
rect 38795 45849 38804 45883
rect 38752 45840 38804 45849
rect 40040 45840 40092 45892
rect 40776 45840 40828 45892
rect 41696 45908 41748 45960
rect 42892 45976 42944 46028
rect 43904 45976 43956 46028
rect 42708 45951 42760 45960
rect 42708 45917 42717 45951
rect 42717 45917 42751 45951
rect 42751 45917 42760 45951
rect 42708 45908 42760 45917
rect 42800 45951 42852 45960
rect 42800 45917 42809 45951
rect 42809 45917 42843 45951
rect 42843 45917 42852 45951
rect 42800 45908 42852 45917
rect 42984 45908 43036 45960
rect 43628 45908 43680 45960
rect 44180 45951 44232 45960
rect 44180 45917 44189 45951
rect 44189 45917 44223 45951
rect 44223 45917 44232 45951
rect 44180 45908 44232 45917
rect 44456 45908 44508 45960
rect 44916 45908 44968 45960
rect 35532 45772 35584 45824
rect 36268 45815 36320 45824
rect 36268 45781 36277 45815
rect 36277 45781 36311 45815
rect 36311 45781 36320 45815
rect 36268 45772 36320 45781
rect 36636 45772 36688 45824
rect 37740 45772 37792 45824
rect 37924 45772 37976 45824
rect 39856 45815 39908 45824
rect 39856 45781 39865 45815
rect 39865 45781 39899 45815
rect 39899 45781 39908 45815
rect 39856 45772 39908 45781
rect 40500 45772 40552 45824
rect 42248 45840 42300 45892
rect 43352 45840 43404 45892
rect 44548 45840 44600 45892
rect 50160 45908 50212 45960
rect 50988 45951 51040 45960
rect 50988 45917 50997 45951
rect 50997 45917 51031 45951
rect 51031 45917 51040 45951
rect 50988 45908 51040 45917
rect 51264 45951 51316 45960
rect 51264 45917 51273 45951
rect 51273 45917 51307 45951
rect 51307 45917 51316 45951
rect 51264 45908 51316 45917
rect 51816 45908 51868 45960
rect 56876 45908 56928 45960
rect 57428 45908 57480 45960
rect 57796 45951 57848 45960
rect 57796 45917 57805 45951
rect 57805 45917 57839 45951
rect 57839 45917 57848 45951
rect 57796 45908 57848 45917
rect 46296 45840 46348 45892
rect 47124 45840 47176 45892
rect 47584 45883 47636 45892
rect 47584 45849 47593 45883
rect 47593 45849 47627 45883
rect 47627 45849 47636 45883
rect 47584 45840 47636 45849
rect 52092 45840 52144 45892
rect 41696 45772 41748 45824
rect 42156 45815 42208 45824
rect 42156 45781 42165 45815
rect 42165 45781 42199 45815
rect 42199 45781 42208 45815
rect 42156 45772 42208 45781
rect 43076 45772 43128 45824
rect 45008 45772 45060 45824
rect 45652 45772 45704 45824
rect 47216 45772 47268 45824
rect 47952 45772 48004 45824
rect 50712 45772 50764 45824
rect 57060 45815 57112 45824
rect 57060 45781 57069 45815
rect 57069 45781 57103 45815
rect 57103 45781 57112 45815
rect 57060 45772 57112 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 20444 45568 20496 45620
rect 2044 45500 2096 45552
rect 22652 45543 22704 45552
rect 18788 45432 18840 45484
rect 20260 45432 20312 45484
rect 20536 45432 20588 45484
rect 20168 45296 20220 45348
rect 20352 45228 20404 45280
rect 22100 45432 22152 45484
rect 22652 45509 22686 45543
rect 22686 45509 22704 45543
rect 22652 45500 22704 45509
rect 25136 45543 25188 45552
rect 25136 45509 25145 45543
rect 25145 45509 25179 45543
rect 25179 45509 25188 45543
rect 25136 45500 25188 45509
rect 25596 45500 25648 45552
rect 33784 45568 33836 45620
rect 22376 45407 22428 45416
rect 22376 45373 22385 45407
rect 22385 45373 22419 45407
rect 22419 45373 22428 45407
rect 22376 45364 22428 45373
rect 25688 45432 25740 45484
rect 28448 45500 28500 45552
rect 30012 45500 30064 45552
rect 33140 45500 33192 45552
rect 37924 45568 37976 45620
rect 38752 45568 38804 45620
rect 39856 45568 39908 45620
rect 28264 45475 28316 45484
rect 28264 45441 28273 45475
rect 28273 45441 28307 45475
rect 28307 45441 28316 45475
rect 28264 45432 28316 45441
rect 34888 45432 34940 45484
rect 39948 45500 40000 45552
rect 40040 45500 40092 45552
rect 24216 45407 24268 45416
rect 24216 45373 24225 45407
rect 24225 45373 24259 45407
rect 24259 45373 24268 45407
rect 29000 45407 29052 45416
rect 24216 45364 24268 45373
rect 25136 45296 25188 45348
rect 29000 45373 29009 45407
rect 29009 45373 29043 45407
rect 29043 45373 29052 45407
rect 29000 45364 29052 45373
rect 31024 45364 31076 45416
rect 32036 45296 32088 45348
rect 24676 45271 24728 45280
rect 24676 45237 24685 45271
rect 24685 45237 24719 45271
rect 24719 45237 24728 45271
rect 24676 45228 24728 45237
rect 24768 45228 24820 45280
rect 26056 45271 26108 45280
rect 26056 45237 26065 45271
rect 26065 45237 26099 45271
rect 26099 45237 26108 45271
rect 26056 45228 26108 45237
rect 34612 45364 34664 45416
rect 33416 45228 33468 45280
rect 33692 45228 33744 45280
rect 35624 45432 35676 45484
rect 36452 45475 36504 45484
rect 36452 45441 36461 45475
rect 36461 45441 36495 45475
rect 36495 45441 36504 45475
rect 36452 45432 36504 45441
rect 36636 45475 36688 45484
rect 36636 45441 36645 45475
rect 36645 45441 36679 45475
rect 36679 45441 36688 45475
rect 36636 45432 36688 45441
rect 36728 45475 36780 45484
rect 36728 45441 36737 45475
rect 36737 45441 36771 45475
rect 36771 45441 36780 45475
rect 36728 45432 36780 45441
rect 37740 45475 37792 45484
rect 37740 45441 37749 45475
rect 37749 45441 37783 45475
rect 37783 45441 37792 45475
rect 37740 45432 37792 45441
rect 38292 45432 38344 45484
rect 38568 45475 38620 45484
rect 38568 45441 38577 45475
rect 38577 45441 38611 45475
rect 38611 45441 38620 45475
rect 38568 45432 38620 45441
rect 39764 45432 39816 45484
rect 40500 45475 40552 45484
rect 40500 45441 40509 45475
rect 40509 45441 40543 45475
rect 40543 45441 40552 45475
rect 40500 45432 40552 45441
rect 35624 45296 35676 45348
rect 39120 45364 39172 45416
rect 37924 45296 37976 45348
rect 38016 45296 38068 45348
rect 35440 45228 35492 45280
rect 35716 45271 35768 45280
rect 35716 45237 35725 45271
rect 35725 45237 35759 45271
rect 35759 45237 35768 45271
rect 35716 45228 35768 45237
rect 35992 45228 36044 45280
rect 36452 45271 36504 45280
rect 36452 45237 36461 45271
rect 36461 45237 36495 45271
rect 36495 45237 36504 45271
rect 36452 45228 36504 45237
rect 37004 45228 37056 45280
rect 38200 45228 38252 45280
rect 38660 45228 38712 45280
rect 40500 45296 40552 45348
rect 40776 45296 40828 45348
rect 41236 45432 41288 45484
rect 42064 45568 42116 45620
rect 42800 45500 42852 45552
rect 40960 45364 41012 45416
rect 41604 45407 41656 45416
rect 41604 45373 41613 45407
rect 41613 45373 41647 45407
rect 41647 45373 41656 45407
rect 41604 45364 41656 45373
rect 41880 45364 41932 45416
rect 42892 45432 42944 45484
rect 43444 45568 43496 45620
rect 43168 45500 43220 45552
rect 45836 45500 45888 45552
rect 48780 45500 48832 45552
rect 49608 45500 49660 45552
rect 45928 45475 45980 45484
rect 45928 45441 45937 45475
rect 45937 45441 45971 45475
rect 45971 45441 45980 45475
rect 45928 45432 45980 45441
rect 46480 45432 46532 45484
rect 47124 45432 47176 45484
rect 43076 45364 43128 45416
rect 46848 45364 46900 45416
rect 47768 45432 47820 45484
rect 48228 45432 48280 45484
rect 48964 45475 49016 45484
rect 48964 45441 48973 45475
rect 48973 45441 49007 45475
rect 49007 45441 49016 45475
rect 48964 45432 49016 45441
rect 49700 45432 49752 45484
rect 51448 45475 51500 45484
rect 51448 45441 51457 45475
rect 51457 45441 51491 45475
rect 51491 45441 51500 45475
rect 51448 45432 51500 45441
rect 55864 45432 55916 45484
rect 56048 45475 56100 45484
rect 56048 45441 56057 45475
rect 56057 45441 56091 45475
rect 56091 45441 56100 45475
rect 56048 45432 56100 45441
rect 47676 45407 47728 45416
rect 47676 45373 47685 45407
rect 47685 45373 47719 45407
rect 47719 45373 47728 45407
rect 47676 45364 47728 45373
rect 48136 45364 48188 45416
rect 51356 45364 51408 45416
rect 51816 45407 51868 45416
rect 47216 45296 47268 45348
rect 48228 45296 48280 45348
rect 49056 45339 49108 45348
rect 49056 45305 49065 45339
rect 49065 45305 49099 45339
rect 49099 45305 49108 45339
rect 49056 45296 49108 45305
rect 51816 45373 51825 45407
rect 51825 45373 51859 45407
rect 51859 45373 51868 45407
rect 51816 45364 51868 45373
rect 52000 45296 52052 45348
rect 42432 45228 42484 45280
rect 45376 45228 45428 45280
rect 45744 45271 45796 45280
rect 45744 45237 45753 45271
rect 45753 45237 45787 45271
rect 45787 45237 45796 45271
rect 45744 45228 45796 45237
rect 47492 45228 47544 45280
rect 47584 45271 47636 45280
rect 47584 45237 47593 45271
rect 47593 45237 47627 45271
rect 47627 45237 47636 45271
rect 47584 45228 47636 45237
rect 52736 45228 52788 45280
rect 55864 45228 55916 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19340 45024 19392 45076
rect 20168 45067 20220 45076
rect 20168 45033 20177 45067
rect 20177 45033 20211 45067
rect 20211 45033 20220 45067
rect 20168 45024 20220 45033
rect 20628 45024 20680 45076
rect 24860 45024 24912 45076
rect 26056 45024 26108 45076
rect 27712 45024 27764 45076
rect 3424 44956 3476 45008
rect 29000 44956 29052 45008
rect 29276 44956 29328 45008
rect 20444 44888 20496 44940
rect 31024 45024 31076 45076
rect 35440 45024 35492 45076
rect 37188 45024 37240 45076
rect 38016 45024 38068 45076
rect 38384 45067 38436 45076
rect 38384 45033 38393 45067
rect 38393 45033 38427 45067
rect 38427 45033 38436 45067
rect 38384 45024 38436 45033
rect 39120 45067 39172 45076
rect 39120 45033 39129 45067
rect 39129 45033 39163 45067
rect 39163 45033 39172 45067
rect 39120 45024 39172 45033
rect 40960 45024 41012 45076
rect 41328 45024 41380 45076
rect 43444 45024 43496 45076
rect 46572 45067 46624 45076
rect 46572 45033 46581 45067
rect 46581 45033 46615 45067
rect 46615 45033 46624 45067
rect 46572 45024 46624 45033
rect 47124 45024 47176 45076
rect 47676 45024 47728 45076
rect 48228 45024 48280 45076
rect 49516 45024 49568 45076
rect 49700 45024 49752 45076
rect 50712 45024 50764 45076
rect 51356 45024 51408 45076
rect 19432 44863 19484 44872
rect 19432 44829 19441 44863
rect 19441 44829 19475 44863
rect 19475 44829 19484 44863
rect 19432 44820 19484 44829
rect 20536 44820 20588 44872
rect 24676 44863 24728 44872
rect 24676 44829 24685 44863
rect 24685 44829 24719 44863
rect 24719 44829 24728 44863
rect 24676 44820 24728 44829
rect 24768 44863 24820 44872
rect 24768 44829 24777 44863
rect 24777 44829 24811 44863
rect 24811 44829 24820 44863
rect 25044 44863 25096 44872
rect 24768 44820 24820 44829
rect 25044 44829 25053 44863
rect 25053 44829 25087 44863
rect 25087 44829 25096 44863
rect 25044 44820 25096 44829
rect 25596 44863 25648 44872
rect 25596 44829 25605 44863
rect 25605 44829 25639 44863
rect 25639 44829 25648 44863
rect 25596 44820 25648 44829
rect 25688 44863 25740 44872
rect 25688 44829 25697 44863
rect 25697 44829 25731 44863
rect 25731 44829 25740 44863
rect 32036 44888 32088 44940
rect 25688 44820 25740 44829
rect 28264 44820 28316 44872
rect 29092 44820 29144 44872
rect 30288 44820 30340 44872
rect 20260 44752 20312 44804
rect 28816 44795 28868 44804
rect 28816 44761 28825 44795
rect 28825 44761 28859 44795
rect 28859 44761 28868 44795
rect 32220 44820 32272 44872
rect 32404 44820 32456 44872
rect 32956 44863 33008 44872
rect 32956 44829 32965 44863
rect 32965 44829 32999 44863
rect 32999 44829 33008 44863
rect 32956 44820 33008 44829
rect 34612 44888 34664 44940
rect 41604 44956 41656 45008
rect 49424 44956 49476 45008
rect 55496 44999 55548 45008
rect 55496 44965 55505 44999
rect 55505 44965 55539 44999
rect 55539 44965 55548 44999
rect 55496 44956 55548 44965
rect 37740 44888 37792 44940
rect 37924 44888 37976 44940
rect 28816 44752 28868 44761
rect 33508 44820 33560 44872
rect 35716 44820 35768 44872
rect 37556 44863 37608 44872
rect 37556 44829 37565 44863
rect 37565 44829 37599 44863
rect 37599 44829 37608 44863
rect 37556 44820 37608 44829
rect 37832 44820 37884 44872
rect 38200 44820 38252 44872
rect 38384 44863 38436 44872
rect 38384 44829 38393 44863
rect 38393 44829 38427 44863
rect 38427 44829 38436 44863
rect 38384 44820 38436 44829
rect 38660 44820 38712 44872
rect 39304 44863 39356 44872
rect 39304 44829 39313 44863
rect 39313 44829 39347 44863
rect 39347 44829 39356 44863
rect 39304 44820 39356 44829
rect 40132 44888 40184 44940
rect 39672 44820 39724 44872
rect 39856 44820 39908 44872
rect 41052 44820 41104 44872
rect 49056 44888 49108 44940
rect 49332 44888 49384 44940
rect 49516 44888 49568 44940
rect 42432 44863 42484 44872
rect 42432 44829 42441 44863
rect 42441 44829 42475 44863
rect 42475 44829 42484 44863
rect 42432 44820 42484 44829
rect 24216 44684 24268 44736
rect 32956 44684 33008 44736
rect 34336 44684 34388 44736
rect 35624 44684 35676 44736
rect 38476 44752 38528 44804
rect 40592 44795 40644 44804
rect 40592 44761 40601 44795
rect 40601 44761 40635 44795
rect 40635 44761 40644 44795
rect 40592 44752 40644 44761
rect 42248 44752 42300 44804
rect 44088 44820 44140 44872
rect 46480 44863 46532 44872
rect 46480 44829 46489 44863
rect 46489 44829 46523 44863
rect 46523 44829 46532 44863
rect 46480 44820 46532 44829
rect 47032 44820 47084 44872
rect 48228 44820 48280 44872
rect 49424 44863 49476 44872
rect 49424 44829 49433 44863
rect 49433 44829 49467 44863
rect 49467 44829 49476 44863
rect 49424 44820 49476 44829
rect 52644 44888 52696 44940
rect 52092 44863 52144 44872
rect 42892 44795 42944 44804
rect 42892 44761 42901 44795
rect 42901 44761 42935 44795
rect 42935 44761 42944 44795
rect 42892 44752 42944 44761
rect 42984 44752 43036 44804
rect 43168 44752 43220 44804
rect 44180 44752 44232 44804
rect 52092 44829 52101 44863
rect 52101 44829 52135 44863
rect 52135 44829 52144 44863
rect 52092 44820 52144 44829
rect 52736 44863 52788 44872
rect 52736 44829 52745 44863
rect 52745 44829 52779 44863
rect 52779 44829 52788 44863
rect 52736 44820 52788 44829
rect 53840 44888 53892 44940
rect 53656 44863 53708 44872
rect 53656 44829 53665 44863
rect 53665 44829 53699 44863
rect 53699 44829 53708 44863
rect 53656 44820 53708 44829
rect 56048 44888 56100 44940
rect 57796 44956 57848 45008
rect 57060 44888 57112 44940
rect 57888 44931 57940 44940
rect 57888 44897 57897 44931
rect 57897 44897 57931 44931
rect 57931 44897 57940 44931
rect 57888 44888 57940 44897
rect 55864 44863 55916 44872
rect 55864 44829 55873 44863
rect 55873 44829 55907 44863
rect 55907 44829 55916 44863
rect 55864 44820 55916 44829
rect 55772 44752 55824 44804
rect 42340 44727 42392 44736
rect 42340 44693 42349 44727
rect 42349 44693 42383 44727
rect 42383 44693 42392 44727
rect 42340 44684 42392 44693
rect 42524 44684 42576 44736
rect 44364 44684 44416 44736
rect 45560 44727 45612 44736
rect 45560 44693 45569 44727
rect 45569 44693 45603 44727
rect 45603 44693 45612 44727
rect 45560 44684 45612 44693
rect 49700 44684 49752 44736
rect 50896 44727 50948 44736
rect 50896 44693 50905 44727
rect 50905 44693 50939 44727
rect 50939 44693 50948 44727
rect 50896 44684 50948 44693
rect 52920 44727 52972 44736
rect 52920 44693 52929 44727
rect 52929 44693 52963 44727
rect 52963 44693 52972 44727
rect 52920 44684 52972 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 19984 44480 20036 44532
rect 24768 44480 24820 44532
rect 38568 44480 38620 44532
rect 39856 44523 39908 44532
rect 39856 44489 39865 44523
rect 39865 44489 39899 44523
rect 39899 44489 39908 44523
rect 39856 44480 39908 44489
rect 40868 44480 40920 44532
rect 41788 44480 41840 44532
rect 2044 44412 2096 44464
rect 2688 44412 2740 44464
rect 20076 44344 20128 44396
rect 27620 44412 27672 44464
rect 24860 44344 24912 44396
rect 25044 44387 25096 44396
rect 25044 44353 25053 44387
rect 25053 44353 25087 44387
rect 25087 44353 25096 44387
rect 25044 44344 25096 44353
rect 31024 44412 31076 44464
rect 32036 44412 32088 44464
rect 29460 44344 29512 44396
rect 32404 44387 32456 44396
rect 32404 44353 32413 44387
rect 32413 44353 32447 44387
rect 32447 44353 32456 44387
rect 32404 44344 32456 44353
rect 37832 44412 37884 44464
rect 39120 44412 39172 44464
rect 40592 44412 40644 44464
rect 32772 44387 32824 44396
rect 32772 44353 32781 44387
rect 32781 44353 32815 44387
rect 32815 44353 32824 44387
rect 32772 44344 32824 44353
rect 33508 44387 33560 44396
rect 33508 44353 33517 44387
rect 33517 44353 33551 44387
rect 33551 44353 33560 44387
rect 33508 44344 33560 44353
rect 35532 44344 35584 44396
rect 35808 44387 35860 44396
rect 35808 44353 35817 44387
rect 35817 44353 35851 44387
rect 35851 44353 35860 44387
rect 35992 44387 36044 44396
rect 35808 44344 35860 44353
rect 35992 44353 36001 44387
rect 36001 44353 36035 44387
rect 36035 44353 36044 44387
rect 35992 44344 36044 44353
rect 39304 44344 39356 44396
rect 41144 44344 41196 44396
rect 41328 44387 41380 44396
rect 41328 44353 41337 44387
rect 41337 44353 41371 44387
rect 41371 44353 41380 44387
rect 41328 44344 41380 44353
rect 41880 44344 41932 44396
rect 42984 44480 43036 44532
rect 43444 44480 43496 44532
rect 44180 44480 44232 44532
rect 44364 44412 44416 44464
rect 47860 44480 47912 44532
rect 48228 44523 48280 44532
rect 48228 44489 48237 44523
rect 48237 44489 48271 44523
rect 48271 44489 48280 44523
rect 48228 44480 48280 44489
rect 48964 44480 49016 44532
rect 50896 44480 50948 44532
rect 52920 44480 52972 44532
rect 53656 44523 53708 44532
rect 53656 44489 53665 44523
rect 53665 44489 53699 44523
rect 53699 44489 53708 44523
rect 53656 44480 53708 44489
rect 24676 44208 24728 44260
rect 32404 44208 32456 44260
rect 2964 44140 3016 44192
rect 3424 44140 3476 44192
rect 24400 44140 24452 44192
rect 30196 44140 30248 44192
rect 32128 44183 32180 44192
rect 32128 44149 32137 44183
rect 32137 44149 32171 44183
rect 32171 44149 32180 44183
rect 32128 44140 32180 44149
rect 34520 44140 34572 44192
rect 38384 44276 38436 44328
rect 42892 44387 42944 44396
rect 42892 44353 42901 44387
rect 42901 44353 42935 44387
rect 42935 44353 42944 44387
rect 42892 44344 42944 44353
rect 43168 44344 43220 44396
rect 43904 44344 43956 44396
rect 44824 44387 44876 44396
rect 44824 44353 44833 44387
rect 44833 44353 44867 44387
rect 44867 44353 44876 44387
rect 44824 44344 44876 44353
rect 45468 44344 45520 44396
rect 47308 44412 47360 44464
rect 46664 44387 46716 44396
rect 46664 44353 46673 44387
rect 46673 44353 46707 44387
rect 46707 44353 46716 44387
rect 46664 44344 46716 44353
rect 43260 44276 43312 44328
rect 43536 44319 43588 44328
rect 43536 44285 43545 44319
rect 43545 44285 43579 44319
rect 43579 44285 43588 44319
rect 43536 44276 43588 44285
rect 43720 44319 43772 44328
rect 43720 44285 43729 44319
rect 43729 44285 43763 44319
rect 43763 44285 43772 44319
rect 43720 44276 43772 44285
rect 38292 44208 38344 44260
rect 41236 44208 41288 44260
rect 41972 44208 42024 44260
rect 42708 44208 42760 44260
rect 45836 44208 45888 44260
rect 46572 44319 46624 44328
rect 46572 44285 46582 44319
rect 46582 44285 46616 44319
rect 46616 44285 46624 44319
rect 48320 44344 48372 44396
rect 48780 44344 48832 44396
rect 49424 44412 49476 44464
rect 50988 44455 51040 44464
rect 50988 44421 50997 44455
rect 50997 44421 51031 44455
rect 51031 44421 51040 44455
rect 50988 44412 51040 44421
rect 51448 44412 51500 44464
rect 49332 44387 49384 44396
rect 49332 44353 49341 44387
rect 49341 44353 49375 44387
rect 49375 44353 49384 44387
rect 49332 44344 49384 44353
rect 50068 44387 50120 44396
rect 50068 44353 50077 44387
rect 50077 44353 50111 44387
rect 50111 44353 50120 44387
rect 50068 44344 50120 44353
rect 46572 44276 46624 44285
rect 48228 44276 48280 44328
rect 50896 44276 50948 44328
rect 52092 44344 52144 44396
rect 52644 44276 52696 44328
rect 47124 44208 47176 44260
rect 52092 44208 52144 44260
rect 53840 44276 53892 44328
rect 55128 44412 55180 44464
rect 56324 44412 56376 44464
rect 55404 44344 55456 44396
rect 56508 44387 56560 44396
rect 56508 44353 56517 44387
rect 56517 44353 56551 44387
rect 56551 44353 56560 44387
rect 56508 44344 56560 44353
rect 56968 44344 57020 44396
rect 55312 44276 55364 44328
rect 55772 44276 55824 44328
rect 39672 44183 39724 44192
rect 39672 44149 39681 44183
rect 39681 44149 39715 44183
rect 39715 44149 39724 44183
rect 39672 44140 39724 44149
rect 42800 44140 42852 44192
rect 46112 44140 46164 44192
rect 47676 44140 47728 44192
rect 53104 44183 53156 44192
rect 53104 44149 53113 44183
rect 53113 44149 53147 44183
rect 53147 44149 53156 44183
rect 53104 44140 53156 44149
rect 54484 44183 54536 44192
rect 54484 44149 54493 44183
rect 54493 44149 54527 44183
rect 54527 44149 54536 44183
rect 54484 44140 54536 44149
rect 56600 44140 56652 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 29460 43936 29512 43988
rect 35532 43936 35584 43988
rect 37556 43936 37608 43988
rect 38936 43936 38988 43988
rect 43720 43936 43772 43988
rect 44824 43936 44876 43988
rect 32772 43868 32824 43920
rect 39028 43868 39080 43920
rect 39120 43868 39172 43920
rect 39764 43868 39816 43920
rect 29092 43800 29144 43852
rect 31024 43800 31076 43852
rect 40316 43843 40368 43852
rect 40316 43809 40325 43843
rect 40325 43809 40359 43843
rect 40359 43809 40368 43843
rect 40316 43800 40368 43809
rect 32128 43732 32180 43784
rect 35900 43732 35952 43784
rect 29092 43664 29144 43716
rect 32404 43596 32456 43648
rect 34612 43596 34664 43648
rect 35992 43596 36044 43648
rect 38108 43775 38160 43784
rect 38108 43741 38117 43775
rect 38117 43741 38151 43775
rect 38151 43741 38160 43775
rect 38752 43775 38804 43784
rect 38108 43732 38160 43741
rect 38752 43741 38761 43775
rect 38761 43741 38795 43775
rect 38795 43741 38804 43775
rect 38752 43732 38804 43741
rect 38936 43775 38988 43784
rect 38936 43741 38945 43775
rect 38945 43741 38979 43775
rect 38979 43741 38988 43775
rect 38936 43732 38988 43741
rect 38292 43664 38344 43716
rect 38384 43664 38436 43716
rect 39764 43732 39816 43784
rect 40040 43775 40092 43784
rect 40040 43741 40049 43775
rect 40049 43741 40083 43775
rect 40083 43741 40092 43775
rect 40040 43732 40092 43741
rect 40684 43732 40736 43784
rect 41144 43732 41196 43784
rect 41972 43800 42024 43852
rect 42156 43868 42208 43920
rect 45560 43868 45612 43920
rect 46020 43936 46072 43988
rect 46848 43868 46900 43920
rect 49332 43868 49384 43920
rect 50068 43936 50120 43988
rect 52644 43979 52696 43988
rect 52644 43945 52653 43979
rect 52653 43945 52687 43979
rect 52687 43945 52696 43979
rect 52644 43936 52696 43945
rect 53840 43979 53892 43988
rect 53840 43945 53849 43979
rect 53849 43945 53883 43979
rect 53883 43945 53892 43979
rect 53840 43936 53892 43945
rect 55128 43936 55180 43988
rect 57152 43936 57204 43988
rect 41052 43664 41104 43716
rect 40960 43596 41012 43648
rect 41328 43596 41380 43648
rect 42432 43732 42484 43784
rect 44916 43800 44968 43852
rect 45192 43843 45244 43852
rect 45192 43809 45201 43843
rect 45201 43809 45235 43843
rect 45235 43809 45244 43843
rect 45192 43800 45244 43809
rect 45652 43800 45704 43852
rect 45744 43800 45796 43852
rect 46756 43843 46808 43852
rect 46756 43809 46765 43843
rect 46765 43809 46799 43843
rect 46799 43809 46808 43843
rect 46756 43800 46808 43809
rect 44180 43775 44232 43784
rect 44180 43741 44189 43775
rect 44189 43741 44223 43775
rect 44223 43741 44232 43775
rect 44180 43732 44232 43741
rect 42800 43707 42852 43716
rect 42800 43673 42809 43707
rect 42809 43673 42843 43707
rect 42843 43673 42852 43707
rect 42800 43664 42852 43673
rect 42984 43664 43036 43716
rect 44916 43664 44968 43716
rect 41696 43596 41748 43648
rect 42616 43596 42668 43648
rect 42892 43639 42944 43648
rect 42892 43605 42901 43639
rect 42901 43605 42935 43639
rect 42935 43605 42944 43639
rect 42892 43596 42944 43605
rect 43996 43596 44048 43648
rect 49608 43800 49660 43852
rect 45376 43664 45428 43716
rect 45652 43707 45704 43716
rect 45652 43673 45661 43707
rect 45661 43673 45695 43707
rect 45695 43673 45704 43707
rect 46480 43732 46532 43784
rect 47584 43732 47636 43784
rect 48136 43732 48188 43784
rect 48596 43732 48648 43784
rect 50068 43732 50120 43784
rect 50988 43800 51040 43852
rect 50620 43732 50672 43784
rect 50804 43775 50856 43784
rect 50804 43741 50813 43775
rect 50813 43741 50847 43775
rect 50847 43741 50856 43775
rect 52276 43775 52328 43784
rect 50804 43732 50856 43741
rect 52276 43741 52285 43775
rect 52285 43741 52319 43775
rect 52319 43741 52328 43775
rect 52276 43732 52328 43741
rect 52920 43732 52972 43784
rect 53840 43732 53892 43784
rect 54300 43732 54352 43784
rect 56600 43800 56652 43852
rect 57888 43843 57940 43852
rect 57888 43809 57897 43843
rect 57897 43809 57931 43843
rect 57931 43809 57940 43843
rect 57888 43800 57940 43809
rect 54484 43732 54536 43784
rect 55312 43707 55364 43716
rect 45652 43664 45704 43673
rect 46204 43596 46256 43648
rect 55312 43673 55321 43707
rect 55321 43673 55355 43707
rect 55355 43673 55364 43707
rect 55312 43664 55364 43673
rect 55956 43664 56008 43716
rect 47860 43596 47912 43648
rect 50620 43596 50672 43648
rect 54760 43639 54812 43648
rect 54760 43605 54769 43639
rect 54769 43605 54803 43639
rect 54803 43605 54812 43639
rect 54760 43596 54812 43605
rect 55404 43596 55456 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 41328 43435 41380 43444
rect 24216 43324 24268 43376
rect 26240 43324 26292 43376
rect 23296 43256 23348 43308
rect 25228 43256 25280 43308
rect 26056 43256 26108 43308
rect 26332 43299 26384 43308
rect 26332 43265 26341 43299
rect 26341 43265 26375 43299
rect 26375 43265 26384 43299
rect 26332 43256 26384 43265
rect 34612 43256 34664 43308
rect 23480 43120 23532 43172
rect 24400 43231 24452 43240
rect 24400 43197 24409 43231
rect 24409 43197 24443 43231
rect 24443 43197 24452 43231
rect 24400 43188 24452 43197
rect 24492 43120 24544 43172
rect 35532 43256 35584 43308
rect 35624 43188 35676 43240
rect 35440 43120 35492 43172
rect 35992 43299 36044 43308
rect 35992 43265 36001 43299
rect 36001 43265 36035 43299
rect 36035 43265 36044 43299
rect 41328 43401 41337 43435
rect 41337 43401 41371 43435
rect 41371 43401 41380 43435
rect 41328 43392 41380 43401
rect 42616 43392 42668 43444
rect 42800 43392 42852 43444
rect 42892 43392 42944 43444
rect 44640 43392 44692 43444
rect 45560 43392 45612 43444
rect 46204 43392 46256 43444
rect 46480 43435 46532 43444
rect 46480 43401 46489 43435
rect 46489 43401 46523 43435
rect 46523 43401 46532 43435
rect 46480 43392 46532 43401
rect 46940 43392 46992 43444
rect 47216 43392 47268 43444
rect 50712 43435 50764 43444
rect 50712 43401 50721 43435
rect 50721 43401 50755 43435
rect 50755 43401 50764 43435
rect 50712 43392 50764 43401
rect 50804 43392 50856 43444
rect 54300 43435 54352 43444
rect 54300 43401 54309 43435
rect 54309 43401 54343 43435
rect 54343 43401 54352 43435
rect 54300 43392 54352 43401
rect 55128 43435 55180 43444
rect 55128 43401 55137 43435
rect 55137 43401 55171 43435
rect 55171 43401 55180 43435
rect 55128 43392 55180 43401
rect 55588 43392 55640 43444
rect 57152 43435 57204 43444
rect 57152 43401 57161 43435
rect 57161 43401 57195 43435
rect 57195 43401 57204 43435
rect 57152 43392 57204 43401
rect 35992 43256 36044 43265
rect 36268 43299 36320 43308
rect 36268 43265 36277 43299
rect 36277 43265 36311 43299
rect 36311 43265 36320 43299
rect 36268 43256 36320 43265
rect 38384 43299 38436 43308
rect 36084 43188 36136 43240
rect 38384 43265 38393 43299
rect 38393 43265 38427 43299
rect 38427 43265 38436 43299
rect 38384 43256 38436 43265
rect 41236 43299 41288 43308
rect 41236 43265 41245 43299
rect 41245 43265 41279 43299
rect 41279 43265 41288 43299
rect 41236 43256 41288 43265
rect 22560 43095 22612 43104
rect 22560 43061 22569 43095
rect 22569 43061 22603 43095
rect 22603 43061 22612 43095
rect 22560 43052 22612 43061
rect 23388 43052 23440 43104
rect 24676 43052 24728 43104
rect 25964 43095 26016 43104
rect 25964 43061 25973 43095
rect 25973 43061 26007 43095
rect 26007 43061 26016 43095
rect 25964 43052 26016 43061
rect 35532 43095 35584 43104
rect 35532 43061 35541 43095
rect 35541 43061 35575 43095
rect 35575 43061 35584 43095
rect 35532 43052 35584 43061
rect 36728 43095 36780 43104
rect 36728 43061 36737 43095
rect 36737 43061 36771 43095
rect 36771 43061 36780 43095
rect 36728 43052 36780 43061
rect 37740 43052 37792 43104
rect 40960 43052 41012 43104
rect 41788 43256 41840 43308
rect 42524 43256 42576 43308
rect 42892 43256 42944 43308
rect 43168 43256 43220 43308
rect 42156 43188 42208 43240
rect 42248 43188 42300 43240
rect 43996 43256 44048 43308
rect 44088 43256 44140 43308
rect 44916 43324 44968 43376
rect 44456 43188 44508 43240
rect 43076 43120 43128 43172
rect 44272 43052 44324 43104
rect 45008 43256 45060 43308
rect 45468 43299 45520 43308
rect 45468 43265 45477 43299
rect 45477 43265 45511 43299
rect 45511 43265 45520 43299
rect 45468 43256 45520 43265
rect 45560 43299 45612 43308
rect 45560 43265 45569 43299
rect 45569 43265 45603 43299
rect 45603 43265 45612 43299
rect 45836 43299 45888 43308
rect 45560 43256 45612 43265
rect 45836 43265 45845 43299
rect 45845 43265 45879 43299
rect 45879 43265 45888 43299
rect 45836 43256 45888 43265
rect 46572 43256 46624 43308
rect 47492 43256 47544 43308
rect 47676 43299 47728 43308
rect 47676 43265 47685 43299
rect 47685 43265 47719 43299
rect 47719 43265 47728 43299
rect 47676 43256 47728 43265
rect 49976 43256 50028 43308
rect 51448 43299 51500 43308
rect 51448 43265 51457 43299
rect 51457 43265 51491 43299
rect 51491 43265 51500 43299
rect 51448 43256 51500 43265
rect 52276 43256 52328 43308
rect 52920 43299 52972 43308
rect 52920 43265 52929 43299
rect 52929 43265 52963 43299
rect 52963 43265 52972 43299
rect 52920 43256 52972 43265
rect 53104 43256 53156 43308
rect 53472 43299 53524 43308
rect 53472 43265 53481 43299
rect 53481 43265 53515 43299
rect 53515 43265 53524 43299
rect 53472 43256 53524 43265
rect 54024 43256 54076 43308
rect 54392 43299 54444 43308
rect 54392 43265 54401 43299
rect 54401 43265 54435 43299
rect 54435 43265 54444 43299
rect 54392 43256 54444 43265
rect 55312 43299 55364 43308
rect 55312 43265 55321 43299
rect 55321 43265 55355 43299
rect 55355 43265 55364 43299
rect 55312 43256 55364 43265
rect 55496 43256 55548 43308
rect 56324 43299 56376 43308
rect 56324 43265 56333 43299
rect 56333 43265 56367 43299
rect 56367 43265 56376 43299
rect 56324 43256 56376 43265
rect 57704 43256 57756 43308
rect 45192 43188 45244 43240
rect 46388 43188 46440 43240
rect 47216 43188 47268 43240
rect 47860 43231 47912 43240
rect 47860 43197 47869 43231
rect 47869 43197 47903 43231
rect 47903 43197 47912 43231
rect 47860 43188 47912 43197
rect 47308 43120 47360 43172
rect 48136 43120 48188 43172
rect 50068 43188 50120 43240
rect 50620 43231 50672 43240
rect 50620 43197 50629 43231
rect 50629 43197 50663 43231
rect 50663 43197 50672 43231
rect 50620 43188 50672 43197
rect 56968 43188 57020 43240
rect 50896 43120 50948 43172
rect 54116 43120 54168 43172
rect 45928 43052 45980 43104
rect 46480 43052 46532 43104
rect 46940 43052 46992 43104
rect 56876 43052 56928 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 21456 42848 21508 42900
rect 23388 42848 23440 42900
rect 33416 42848 33468 42900
rect 37740 42891 37792 42900
rect 37740 42857 37749 42891
rect 37749 42857 37783 42891
rect 37783 42857 37792 42891
rect 37740 42848 37792 42857
rect 40040 42848 40092 42900
rect 41236 42848 41288 42900
rect 22744 42780 22796 42832
rect 23296 42780 23348 42832
rect 23664 42823 23716 42832
rect 23664 42789 23673 42823
rect 23673 42789 23707 42823
rect 23707 42789 23716 42823
rect 23664 42780 23716 42789
rect 24952 42780 25004 42832
rect 35900 42780 35952 42832
rect 41604 42780 41656 42832
rect 41788 42780 41840 42832
rect 20628 42755 20680 42764
rect 20260 42687 20312 42696
rect 20260 42653 20269 42687
rect 20269 42653 20303 42687
rect 20303 42653 20312 42687
rect 20260 42644 20312 42653
rect 20628 42721 20637 42755
rect 20637 42721 20671 42755
rect 20671 42721 20680 42755
rect 20628 42712 20680 42721
rect 21180 42687 21232 42696
rect 21180 42653 21189 42687
rect 21189 42653 21223 42687
rect 21223 42653 21232 42687
rect 21180 42644 21232 42653
rect 23388 42712 23440 42764
rect 30932 42712 30984 42764
rect 31944 42755 31996 42764
rect 22836 42644 22888 42696
rect 23480 42687 23532 42696
rect 23480 42653 23489 42687
rect 23489 42653 23523 42687
rect 23523 42653 23532 42687
rect 23480 42644 23532 42653
rect 23756 42687 23808 42696
rect 23756 42653 23765 42687
rect 23765 42653 23799 42687
rect 23799 42653 23808 42687
rect 23756 42644 23808 42653
rect 24308 42644 24360 42696
rect 21272 42576 21324 42628
rect 24492 42644 24544 42696
rect 24676 42687 24728 42696
rect 24676 42653 24685 42687
rect 24685 42653 24719 42687
rect 24719 42653 24728 42687
rect 24676 42644 24728 42653
rect 28080 42644 28132 42696
rect 29000 42644 29052 42696
rect 30196 42687 30248 42696
rect 30196 42653 30205 42687
rect 30205 42653 30239 42687
rect 30239 42653 30248 42687
rect 30196 42644 30248 42653
rect 31300 42644 31352 42696
rect 31576 42687 31628 42696
rect 31576 42653 31585 42687
rect 31585 42653 31619 42687
rect 31619 42653 31628 42687
rect 31576 42644 31628 42653
rect 31944 42721 31953 42755
rect 31953 42721 31987 42755
rect 31987 42721 31996 42755
rect 31944 42712 31996 42721
rect 32680 42755 32732 42764
rect 32680 42721 32689 42755
rect 32689 42721 32723 42755
rect 32723 42721 32732 42755
rect 32680 42712 32732 42721
rect 37556 42755 37608 42764
rect 37556 42721 37565 42755
rect 37565 42721 37599 42755
rect 37599 42721 37608 42755
rect 37556 42712 37608 42721
rect 38384 42755 38436 42764
rect 38384 42721 38393 42755
rect 38393 42721 38427 42755
rect 38427 42721 38436 42755
rect 38384 42712 38436 42721
rect 42248 42848 42300 42900
rect 42708 42848 42760 42900
rect 45376 42848 45428 42900
rect 46388 42848 46440 42900
rect 46756 42848 46808 42900
rect 49792 42848 49844 42900
rect 51448 42848 51500 42900
rect 52920 42848 52972 42900
rect 55404 42891 55456 42900
rect 55404 42857 55413 42891
rect 55413 42857 55447 42891
rect 55447 42857 55456 42891
rect 55404 42848 55456 42857
rect 44272 42780 44324 42832
rect 54760 42780 54812 42832
rect 42800 42712 42852 42764
rect 44456 42712 44508 42764
rect 34704 42687 34756 42696
rect 34704 42653 34713 42687
rect 34713 42653 34747 42687
rect 34747 42653 34756 42687
rect 34704 42644 34756 42653
rect 36728 42644 36780 42696
rect 25780 42576 25832 42628
rect 24492 42551 24544 42560
rect 24492 42517 24507 42551
rect 24507 42517 24541 42551
rect 24541 42517 24544 42551
rect 24492 42508 24544 42517
rect 27436 42619 27488 42628
rect 27436 42585 27445 42619
rect 27445 42585 27479 42619
rect 27479 42585 27488 42619
rect 27436 42576 27488 42585
rect 29368 42508 29420 42560
rect 29460 42508 29512 42560
rect 32312 42508 32364 42560
rect 32956 42508 33008 42560
rect 36084 42551 36136 42560
rect 36084 42517 36093 42551
rect 36093 42517 36127 42551
rect 36127 42517 36136 42551
rect 36084 42508 36136 42517
rect 38568 42644 38620 42696
rect 41420 42687 41472 42696
rect 41420 42653 41462 42687
rect 41462 42653 41472 42687
rect 41420 42644 41472 42653
rect 42064 42644 42116 42696
rect 44364 42644 44416 42696
rect 45008 42687 45060 42696
rect 45008 42653 45017 42687
rect 45017 42653 45051 42687
rect 45051 42653 45060 42687
rect 45008 42644 45060 42653
rect 45192 42687 45244 42696
rect 45192 42653 45201 42687
rect 45201 42653 45235 42687
rect 45235 42653 45244 42687
rect 45192 42644 45244 42653
rect 38660 42576 38712 42628
rect 39672 42576 39724 42628
rect 43076 42576 43128 42628
rect 41144 42508 41196 42560
rect 42892 42508 42944 42560
rect 45192 42508 45244 42560
rect 45376 42687 45428 42696
rect 45376 42653 45385 42687
rect 45385 42653 45419 42687
rect 45419 42653 45428 42687
rect 45560 42687 45612 42696
rect 45376 42644 45428 42653
rect 45560 42653 45569 42687
rect 45569 42653 45603 42687
rect 45603 42653 45612 42687
rect 45560 42644 45612 42653
rect 46572 42644 46624 42696
rect 47124 42687 47176 42696
rect 47124 42653 47133 42687
rect 47133 42653 47167 42687
rect 47167 42653 47176 42687
rect 47124 42644 47176 42653
rect 47308 42687 47360 42696
rect 47308 42653 47317 42687
rect 47317 42653 47351 42687
rect 47351 42653 47360 42687
rect 47308 42644 47360 42653
rect 48136 42687 48188 42696
rect 48136 42653 48145 42687
rect 48145 42653 48179 42687
rect 48179 42653 48188 42687
rect 48136 42644 48188 42653
rect 48320 42687 48372 42696
rect 48320 42653 48329 42687
rect 48329 42653 48363 42687
rect 48363 42653 48372 42687
rect 48320 42644 48372 42653
rect 49976 42644 50028 42696
rect 53840 42712 53892 42764
rect 56876 42712 56928 42764
rect 57888 42755 57940 42764
rect 57888 42721 57897 42755
rect 57897 42721 57931 42755
rect 57931 42721 57940 42755
rect 57888 42712 57940 42721
rect 46480 42619 46532 42628
rect 46480 42585 46489 42619
rect 46489 42585 46523 42619
rect 46523 42585 46532 42619
rect 46480 42576 46532 42585
rect 50620 42619 50672 42628
rect 50620 42585 50629 42619
rect 50629 42585 50663 42619
rect 50663 42585 50672 42619
rect 50620 42576 50672 42585
rect 50804 42576 50856 42628
rect 53472 42644 53524 42696
rect 55588 42687 55640 42696
rect 55588 42653 55597 42687
rect 55597 42653 55631 42687
rect 55631 42653 55640 42687
rect 55588 42644 55640 42653
rect 53104 42576 53156 42628
rect 54024 42619 54076 42628
rect 54024 42585 54033 42619
rect 54033 42585 54067 42619
rect 54067 42585 54076 42619
rect 54024 42576 54076 42585
rect 48228 42508 48280 42560
rect 51540 42508 51592 42560
rect 54392 42576 54444 42628
rect 55312 42619 55364 42628
rect 55312 42585 55321 42619
rect 55321 42585 55355 42619
rect 55355 42585 55364 42619
rect 55312 42576 55364 42585
rect 55496 42619 55548 42628
rect 55496 42585 55505 42619
rect 55505 42585 55539 42619
rect 55539 42585 55548 42619
rect 55496 42576 55548 42585
rect 58072 42576 58124 42628
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 20260 42304 20312 42356
rect 23480 42304 23532 42356
rect 25228 42347 25280 42356
rect 25228 42313 25237 42347
rect 25237 42313 25271 42347
rect 25271 42313 25280 42347
rect 25228 42304 25280 42313
rect 25780 42347 25832 42356
rect 25780 42313 25789 42347
rect 25789 42313 25823 42347
rect 25823 42313 25832 42347
rect 25780 42304 25832 42313
rect 29552 42347 29604 42356
rect 29552 42313 29561 42347
rect 29561 42313 29595 42347
rect 29595 42313 29604 42347
rect 29552 42304 29604 42313
rect 21180 42236 21232 42288
rect 22376 42236 22428 42288
rect 23388 42236 23440 42288
rect 20168 42168 20220 42220
rect 22008 42211 22060 42220
rect 22008 42177 22017 42211
rect 22017 42177 22051 42211
rect 22051 42177 22060 42211
rect 22008 42168 22060 42177
rect 23940 42168 23992 42220
rect 25964 42211 26016 42220
rect 25964 42177 25973 42211
rect 25973 42177 26007 42211
rect 26007 42177 26016 42211
rect 25964 42168 26016 42177
rect 26240 42211 26292 42220
rect 26240 42177 26249 42211
rect 26249 42177 26283 42211
rect 26283 42177 26292 42211
rect 26240 42168 26292 42177
rect 26332 42168 26384 42220
rect 27436 42168 27488 42220
rect 27528 42211 27580 42220
rect 27528 42177 27537 42211
rect 27537 42177 27571 42211
rect 27571 42177 27580 42211
rect 28264 42211 28316 42220
rect 27528 42168 27580 42177
rect 28264 42177 28273 42211
rect 28273 42177 28307 42211
rect 28307 42177 28316 42211
rect 28264 42168 28316 42177
rect 29828 42168 29880 42220
rect 31392 42211 31444 42220
rect 20628 42100 20680 42152
rect 30472 42100 30524 42152
rect 31392 42177 31401 42211
rect 31401 42177 31435 42211
rect 31435 42177 31444 42211
rect 31392 42168 31444 42177
rect 32680 42304 32732 42356
rect 35624 42347 35676 42356
rect 35624 42313 35633 42347
rect 35633 42313 35667 42347
rect 35667 42313 35676 42347
rect 35624 42304 35676 42313
rect 38936 42304 38988 42356
rect 42064 42304 42116 42356
rect 42800 42347 42852 42356
rect 42800 42313 42809 42347
rect 42809 42313 42843 42347
rect 42843 42313 42852 42347
rect 42800 42304 42852 42313
rect 47124 42304 47176 42356
rect 49240 42304 49292 42356
rect 50068 42347 50120 42356
rect 50068 42313 50077 42347
rect 50077 42313 50111 42347
rect 50111 42313 50120 42347
rect 50068 42304 50120 42313
rect 52276 42304 52328 42356
rect 54024 42304 54076 42356
rect 55588 42304 55640 42356
rect 56968 42347 57020 42356
rect 56968 42313 56977 42347
rect 56977 42313 57011 42347
rect 57011 42313 57020 42347
rect 56968 42304 57020 42313
rect 32404 42279 32456 42288
rect 32404 42245 32413 42279
rect 32413 42245 32447 42279
rect 32447 42245 32456 42279
rect 32404 42236 32456 42245
rect 32496 42211 32548 42220
rect 32496 42177 32505 42211
rect 32505 42177 32539 42211
rect 32539 42177 32548 42211
rect 32496 42168 32548 42177
rect 34704 42236 34756 42288
rect 39304 42279 39356 42288
rect 39304 42245 39313 42279
rect 39313 42245 39347 42279
rect 39347 42245 39356 42279
rect 39304 42236 39356 42245
rect 42432 42279 42484 42288
rect 42432 42245 42441 42279
rect 42441 42245 42475 42279
rect 42475 42245 42484 42279
rect 42432 42236 42484 42245
rect 48596 42279 48648 42288
rect 35532 42168 35584 42220
rect 37832 42168 37884 42220
rect 38200 42168 38252 42220
rect 39120 42211 39172 42220
rect 39120 42177 39129 42211
rect 39129 42177 39163 42211
rect 39163 42177 39172 42211
rect 39120 42168 39172 42177
rect 33508 42100 33560 42152
rect 41144 42168 41196 42220
rect 41696 42100 41748 42152
rect 32036 42032 32088 42084
rect 22284 42007 22336 42016
rect 22284 41973 22293 42007
rect 22293 41973 22327 42007
rect 22327 41973 22336 42007
rect 22284 41964 22336 41973
rect 24584 41964 24636 42016
rect 27712 42007 27764 42016
rect 27712 41973 27721 42007
rect 27721 41973 27755 42007
rect 27755 41973 27764 42007
rect 27712 41964 27764 41973
rect 30380 41964 30432 42016
rect 31208 42007 31260 42016
rect 31208 41973 31217 42007
rect 31217 41973 31251 42007
rect 31251 41973 31260 42007
rect 31208 41964 31260 41973
rect 32404 41964 32456 42016
rect 32772 41964 32824 42016
rect 39672 41964 39724 42016
rect 41880 42211 41932 42220
rect 41880 42177 41889 42211
rect 41889 42177 41923 42211
rect 41923 42177 41932 42211
rect 48596 42245 48605 42279
rect 48605 42245 48639 42279
rect 48639 42245 48648 42279
rect 48596 42236 48648 42245
rect 56508 42236 56560 42288
rect 43260 42211 43312 42220
rect 41880 42168 41932 42177
rect 43260 42177 43269 42211
rect 43269 42177 43303 42211
rect 43303 42177 43312 42211
rect 43260 42168 43312 42177
rect 43444 42211 43496 42220
rect 43444 42177 43453 42211
rect 43453 42177 43487 42211
rect 43487 42177 43496 42211
rect 43444 42168 43496 42177
rect 47768 42211 47820 42220
rect 47768 42177 47777 42211
rect 47777 42177 47811 42211
rect 47811 42177 47820 42211
rect 47768 42168 47820 42177
rect 48504 42211 48556 42220
rect 48504 42177 48513 42211
rect 48513 42177 48547 42211
rect 48547 42177 48556 42211
rect 48504 42168 48556 42177
rect 46480 42100 46532 42152
rect 48872 42168 48924 42220
rect 49976 42211 50028 42220
rect 49976 42177 49985 42211
rect 49985 42177 50019 42211
rect 50019 42177 50028 42211
rect 49976 42168 50028 42177
rect 49792 42100 49844 42152
rect 50804 42168 50856 42220
rect 51540 42168 51592 42220
rect 51908 42211 51960 42220
rect 51908 42177 51917 42211
rect 51917 42177 51951 42211
rect 51951 42177 51960 42211
rect 51908 42168 51960 42177
rect 54116 42211 54168 42220
rect 54116 42177 54125 42211
rect 54125 42177 54159 42211
rect 54159 42177 54168 42211
rect 54116 42168 54168 42177
rect 55128 42168 55180 42220
rect 58072 42211 58124 42220
rect 58072 42177 58081 42211
rect 58081 42177 58115 42211
rect 58115 42177 58124 42211
rect 58072 42168 58124 42177
rect 57336 42100 57388 42152
rect 42432 42032 42484 42084
rect 47308 42032 47360 42084
rect 47860 42032 47912 42084
rect 50160 42032 50212 42084
rect 50804 42032 50856 42084
rect 42708 41964 42760 42016
rect 54116 41964 54168 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 20168 41803 20220 41812
rect 20168 41769 20177 41803
rect 20177 41769 20211 41803
rect 20211 41769 20220 41803
rect 20168 41760 20220 41769
rect 20996 41760 21048 41812
rect 21272 41803 21324 41812
rect 21272 41769 21281 41803
rect 21281 41769 21315 41803
rect 21315 41769 21324 41803
rect 21272 41760 21324 41769
rect 22008 41760 22060 41812
rect 23940 41760 23992 41812
rect 24952 41803 25004 41812
rect 24952 41769 24961 41803
rect 24961 41769 24995 41803
rect 24995 41769 25004 41803
rect 24952 41760 25004 41769
rect 27528 41760 27580 41812
rect 28080 41803 28132 41812
rect 28080 41769 28089 41803
rect 28089 41769 28123 41803
rect 28123 41769 28132 41803
rect 28080 41760 28132 41769
rect 29000 41803 29052 41812
rect 29000 41769 29009 41803
rect 29009 41769 29043 41803
rect 29043 41769 29052 41803
rect 29000 41760 29052 41769
rect 31300 41760 31352 41812
rect 29920 41692 29972 41744
rect 31208 41692 31260 41744
rect 38384 41760 38436 41812
rect 43260 41760 43312 41812
rect 48320 41760 48372 41812
rect 56508 41760 56560 41812
rect 19984 41556 20036 41608
rect 20444 41599 20496 41608
rect 20444 41565 20453 41599
rect 20453 41565 20487 41599
rect 20487 41565 20496 41599
rect 20444 41556 20496 41565
rect 21180 41624 21232 41676
rect 20812 41599 20864 41608
rect 20812 41565 20821 41599
rect 20821 41565 20855 41599
rect 20855 41565 20864 41599
rect 22376 41624 22428 41676
rect 25044 41624 25096 41676
rect 20812 41556 20864 41565
rect 21732 41599 21784 41608
rect 21732 41565 21746 41599
rect 21746 41565 21780 41599
rect 21780 41565 21784 41599
rect 21732 41556 21784 41565
rect 21916 41599 21968 41608
rect 21916 41565 21925 41599
rect 21925 41565 21959 41599
rect 21959 41565 21968 41599
rect 21916 41556 21968 41565
rect 22192 41556 22244 41608
rect 22836 41599 22888 41608
rect 22836 41565 22845 41599
rect 22845 41565 22879 41599
rect 22879 41565 22888 41599
rect 22836 41556 22888 41565
rect 24124 41556 24176 41608
rect 25228 41556 25280 41608
rect 27988 41624 28040 41676
rect 28540 41667 28592 41676
rect 28540 41633 28549 41667
rect 28549 41633 28583 41667
rect 28583 41633 28592 41667
rect 28540 41624 28592 41633
rect 29368 41624 29420 41676
rect 28908 41556 28960 41608
rect 29000 41556 29052 41608
rect 33600 41692 33652 41744
rect 42524 41692 42576 41744
rect 32588 41667 32640 41676
rect 32588 41633 32597 41667
rect 32597 41633 32631 41667
rect 32631 41633 32640 41667
rect 32588 41624 32640 41633
rect 21088 41420 21140 41472
rect 21456 41488 21508 41540
rect 22744 41531 22796 41540
rect 22744 41497 22753 41531
rect 22753 41497 22787 41531
rect 22787 41497 22796 41531
rect 22744 41488 22796 41497
rect 24768 41488 24820 41540
rect 31116 41488 31168 41540
rect 31576 41488 31628 41540
rect 32312 41565 32322 41586
rect 32322 41565 32356 41586
rect 32356 41565 32364 41586
rect 32312 41534 32364 41565
rect 32680 41556 32732 41608
rect 37280 41599 37332 41608
rect 37280 41565 37289 41599
rect 37289 41565 37323 41599
rect 37323 41565 37332 41599
rect 37280 41556 37332 41565
rect 37556 41599 37608 41608
rect 37556 41565 37565 41599
rect 37565 41565 37599 41599
rect 37599 41565 37608 41599
rect 37556 41556 37608 41565
rect 37924 41556 37976 41608
rect 39304 41556 39356 41608
rect 42432 41599 42484 41608
rect 42432 41565 42441 41599
rect 42441 41565 42475 41599
rect 42475 41565 42484 41599
rect 42432 41556 42484 41565
rect 43168 41556 43220 41608
rect 45560 41624 45612 41676
rect 47676 41624 47728 41676
rect 47952 41692 48004 41744
rect 51080 41624 51132 41676
rect 45192 41599 45244 41608
rect 45192 41565 45201 41599
rect 45201 41565 45235 41599
rect 45235 41565 45244 41599
rect 45192 41556 45244 41565
rect 21824 41420 21876 41472
rect 24584 41420 24636 41472
rect 25044 41420 25096 41472
rect 31944 41463 31996 41472
rect 31944 41429 31953 41463
rect 31953 41429 31987 41463
rect 31987 41429 31996 41463
rect 31944 41420 31996 41429
rect 32128 41420 32180 41472
rect 39948 41488 40000 41540
rect 42340 41488 42392 41540
rect 42892 41488 42944 41540
rect 47308 41488 47360 41540
rect 48504 41556 48556 41608
rect 50068 41556 50120 41608
rect 50712 41599 50764 41608
rect 50712 41565 50721 41599
rect 50721 41565 50755 41599
rect 50755 41565 50764 41599
rect 50712 41556 50764 41565
rect 51172 41599 51224 41608
rect 51172 41565 51181 41599
rect 51181 41565 51215 41599
rect 51215 41565 51224 41599
rect 51172 41556 51224 41565
rect 57244 41556 57296 41608
rect 52552 41488 52604 41540
rect 57152 41488 57204 41540
rect 32588 41420 32640 41472
rect 33048 41420 33100 41472
rect 38660 41420 38712 41472
rect 42616 41420 42668 41472
rect 45284 41463 45336 41472
rect 45284 41429 45293 41463
rect 45293 41429 45327 41463
rect 45327 41429 45336 41463
rect 45284 41420 45336 41429
rect 47400 41420 47452 41472
rect 50988 41420 51040 41472
rect 51080 41420 51132 41472
rect 51448 41420 51500 41472
rect 56784 41420 56836 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 22192 41259 22244 41268
rect 22192 41225 22201 41259
rect 22201 41225 22235 41259
rect 22235 41225 22244 41259
rect 22192 41216 22244 41225
rect 24860 41216 24912 41268
rect 27528 41216 27580 41268
rect 30840 41216 30892 41268
rect 33508 41259 33560 41268
rect 33508 41225 33517 41259
rect 33517 41225 33551 41259
rect 33551 41225 33560 41259
rect 33508 41216 33560 41225
rect 33600 41216 33652 41268
rect 38200 41216 38252 41268
rect 39120 41216 39172 41268
rect 22744 41148 22796 41200
rect 29276 41148 29328 41200
rect 32312 41191 32364 41200
rect 23940 41123 23992 41132
rect 23940 41089 23949 41123
rect 23949 41089 23983 41123
rect 23983 41089 23992 41123
rect 23940 41080 23992 41089
rect 24124 41123 24176 41132
rect 24124 41089 24133 41123
rect 24133 41089 24167 41123
rect 24167 41089 24176 41123
rect 24124 41080 24176 41089
rect 24584 41123 24636 41132
rect 24584 41089 24593 41123
rect 24593 41089 24627 41123
rect 24627 41089 24636 41123
rect 24584 41080 24636 41089
rect 29552 41080 29604 41132
rect 29828 41123 29880 41132
rect 20536 41055 20588 41064
rect 20536 41021 20545 41055
rect 20545 41021 20579 41055
rect 20579 41021 20588 41055
rect 20536 41012 20588 41021
rect 20996 41055 21048 41064
rect 20996 41021 21005 41055
rect 21005 41021 21039 41055
rect 21039 41021 21048 41055
rect 20996 41012 21048 41021
rect 19984 40944 20036 40996
rect 23664 41012 23716 41064
rect 24952 41012 25004 41064
rect 26424 41012 26476 41064
rect 27620 41055 27672 41064
rect 27620 41021 27629 41055
rect 27629 41021 27663 41055
rect 27663 41021 27672 41055
rect 27620 41012 27672 41021
rect 29828 41089 29837 41123
rect 29837 41089 29871 41123
rect 29871 41089 29880 41123
rect 29828 41080 29880 41089
rect 30196 41080 30248 41132
rect 30472 41080 30524 41132
rect 31392 41012 31444 41064
rect 24768 40987 24820 40996
rect 24768 40953 24777 40987
rect 24777 40953 24811 40987
rect 24811 40953 24820 40987
rect 24768 40944 24820 40953
rect 29184 40944 29236 40996
rect 30012 40944 30064 40996
rect 30196 40944 30248 40996
rect 24676 40919 24728 40928
rect 24676 40885 24685 40919
rect 24685 40885 24719 40919
rect 24719 40885 24728 40919
rect 24676 40876 24728 40885
rect 28356 40876 28408 40928
rect 30748 40876 30800 40928
rect 32312 41157 32321 41191
rect 32321 41157 32355 41191
rect 32355 41157 32364 41191
rect 32312 41148 32364 41157
rect 35624 41148 35676 41200
rect 39948 41216 40000 41268
rect 41696 41216 41748 41268
rect 43444 41216 43496 41268
rect 49240 41259 49292 41268
rect 32128 41123 32180 41132
rect 32128 41089 32137 41123
rect 32137 41089 32171 41123
rect 32171 41089 32180 41123
rect 32128 41080 32180 41089
rect 32588 41080 32640 41132
rect 33140 41123 33192 41132
rect 33140 41089 33149 41123
rect 33149 41089 33183 41123
rect 33183 41089 33192 41123
rect 33140 41080 33192 41089
rect 33416 41080 33468 41132
rect 34152 41123 34204 41132
rect 34152 41089 34161 41123
rect 34161 41089 34195 41123
rect 34195 41089 34204 41123
rect 34152 41080 34204 41089
rect 37924 41080 37976 41132
rect 38476 41080 38528 41132
rect 31852 40944 31904 40996
rect 37832 41012 37884 41064
rect 40684 41080 40736 41132
rect 41420 41080 41472 41132
rect 40868 41012 40920 41064
rect 41604 41080 41656 41132
rect 41788 41080 41840 41132
rect 42892 41123 42944 41132
rect 42892 41089 42901 41123
rect 42901 41089 42935 41123
rect 42935 41089 42944 41123
rect 42892 41080 42944 41089
rect 42432 41012 42484 41064
rect 45928 41080 45980 41132
rect 46296 41080 46348 41132
rect 47124 41148 47176 41200
rect 49240 41225 49249 41259
rect 49249 41225 49283 41259
rect 49283 41225 49292 41259
rect 49240 41216 49292 41225
rect 49608 41148 49660 41200
rect 51172 41216 51224 41268
rect 51540 41259 51592 41268
rect 51540 41225 51549 41259
rect 51549 41225 51583 41259
rect 51583 41225 51592 41259
rect 51540 41216 51592 41225
rect 55312 41216 55364 41268
rect 57336 41216 57388 41268
rect 51908 41148 51960 41200
rect 56784 41148 56836 41200
rect 57152 41148 57204 41200
rect 47400 41080 47452 41132
rect 41696 40944 41748 40996
rect 47216 41012 47268 41064
rect 48228 41123 48280 41132
rect 48228 41089 48242 41123
rect 48242 41089 48276 41123
rect 48276 41089 48280 41123
rect 48228 41080 48280 41089
rect 49240 41080 49292 41132
rect 50068 41123 50120 41132
rect 50068 41089 50074 41123
rect 50074 41089 50108 41123
rect 50108 41089 50120 41123
rect 50988 41123 51040 41132
rect 50068 41080 50120 41089
rect 50988 41089 50997 41123
rect 50997 41089 51031 41123
rect 51031 41089 51040 41123
rect 50988 41080 51040 41089
rect 48688 41012 48740 41064
rect 50528 41055 50580 41064
rect 49516 40944 49568 40996
rect 50528 41021 50537 41055
rect 50537 41021 50571 41055
rect 50571 41021 50580 41055
rect 50528 41012 50580 41021
rect 51080 40944 51132 40996
rect 52184 41123 52236 41132
rect 52184 41089 52193 41123
rect 52193 41089 52227 41123
rect 52227 41089 52236 41123
rect 52184 41080 52236 41089
rect 56232 41123 56284 41132
rect 56232 41089 56241 41123
rect 56241 41089 56275 41123
rect 56275 41089 56284 41123
rect 56232 41080 56284 41089
rect 57244 41080 57296 41132
rect 52460 41012 52512 41064
rect 52736 40944 52788 40996
rect 38568 40876 38620 40928
rect 46940 40919 46992 40928
rect 46940 40885 46949 40919
rect 46949 40885 46983 40919
rect 46983 40885 46992 40919
rect 46940 40876 46992 40885
rect 47400 40876 47452 40928
rect 49424 40876 49476 40928
rect 51632 40876 51684 40928
rect 57244 40876 57296 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 21088 40715 21140 40724
rect 21088 40681 21097 40715
rect 21097 40681 21131 40715
rect 21131 40681 21140 40715
rect 21088 40672 21140 40681
rect 21732 40672 21784 40724
rect 21824 40715 21876 40724
rect 21824 40681 21833 40715
rect 21833 40681 21867 40715
rect 21867 40681 21876 40715
rect 29920 40715 29972 40724
rect 21824 40672 21876 40681
rect 29920 40681 29929 40715
rect 29929 40681 29963 40715
rect 29963 40681 29972 40715
rect 29920 40672 29972 40681
rect 31300 40715 31352 40724
rect 31300 40681 31309 40715
rect 31309 40681 31343 40715
rect 31343 40681 31352 40715
rect 31300 40672 31352 40681
rect 31760 40672 31812 40724
rect 21916 40604 21968 40656
rect 22652 40604 22704 40656
rect 31392 40604 31444 40656
rect 37280 40672 37332 40724
rect 40776 40672 40828 40724
rect 42708 40672 42760 40724
rect 47952 40672 48004 40724
rect 49516 40715 49568 40724
rect 49516 40681 49525 40715
rect 49525 40681 49559 40715
rect 49559 40681 49568 40715
rect 49516 40672 49568 40681
rect 49608 40672 49660 40724
rect 52460 40672 52512 40724
rect 56232 40672 56284 40724
rect 57244 40715 57296 40724
rect 57244 40681 57253 40715
rect 57253 40681 57287 40715
rect 57287 40681 57296 40715
rect 57244 40672 57296 40681
rect 33876 40604 33928 40656
rect 34888 40604 34940 40656
rect 22284 40536 22336 40588
rect 23664 40536 23716 40588
rect 24492 40536 24544 40588
rect 27988 40536 28040 40588
rect 30104 40536 30156 40588
rect 21916 40511 21968 40520
rect 21916 40477 21925 40511
rect 21925 40477 21959 40511
rect 21959 40477 21968 40511
rect 21916 40468 21968 40477
rect 24308 40468 24360 40520
rect 25412 40468 25464 40520
rect 28356 40511 28408 40520
rect 22192 40400 22244 40452
rect 22744 40400 22796 40452
rect 23756 40400 23808 40452
rect 25504 40443 25556 40452
rect 25504 40409 25513 40443
rect 25513 40409 25547 40443
rect 25547 40409 25556 40443
rect 25504 40400 25556 40409
rect 28356 40477 28365 40511
rect 28365 40477 28399 40511
rect 28399 40477 28408 40511
rect 28356 40468 28408 40477
rect 31760 40536 31812 40588
rect 31668 40468 31720 40520
rect 33140 40536 33192 40588
rect 32496 40468 32548 40520
rect 32680 40468 32732 40520
rect 33600 40468 33652 40520
rect 37832 40536 37884 40588
rect 37924 40536 37976 40588
rect 40224 40604 40276 40656
rect 31116 40443 31168 40452
rect 31116 40409 31125 40443
rect 31125 40409 31159 40443
rect 31159 40409 31168 40443
rect 31116 40400 31168 40409
rect 32588 40400 32640 40452
rect 34980 40400 35032 40452
rect 37188 40511 37240 40520
rect 37188 40477 37197 40511
rect 37197 40477 37231 40511
rect 37231 40477 37240 40511
rect 38568 40511 38620 40520
rect 37188 40468 37240 40477
rect 38568 40477 38577 40511
rect 38577 40477 38611 40511
rect 38611 40477 38620 40511
rect 38568 40468 38620 40477
rect 39948 40536 40000 40588
rect 40868 40536 40920 40588
rect 39120 40511 39172 40520
rect 39120 40477 39129 40511
rect 39129 40477 39163 40511
rect 39163 40477 39172 40511
rect 39120 40468 39172 40477
rect 22284 40332 22336 40384
rect 26240 40332 26292 40384
rect 27896 40332 27948 40384
rect 30380 40332 30432 40384
rect 30472 40332 30524 40384
rect 33140 40332 33192 40384
rect 33876 40332 33928 40384
rect 34796 40332 34848 40384
rect 37188 40332 37240 40384
rect 38752 40332 38804 40384
rect 39120 40332 39172 40384
rect 39488 40332 39540 40384
rect 41604 40468 41656 40520
rect 41696 40511 41748 40520
rect 41696 40477 41717 40511
rect 41717 40477 41748 40511
rect 43168 40536 43220 40588
rect 46848 40536 46900 40588
rect 42156 40511 42208 40520
rect 41696 40468 41748 40477
rect 42156 40477 42165 40511
rect 42165 40477 42199 40511
rect 42199 40477 42208 40511
rect 42156 40468 42208 40477
rect 42248 40468 42300 40520
rect 42892 40511 42944 40520
rect 42892 40477 42901 40511
rect 42901 40477 42935 40511
rect 42935 40477 42944 40511
rect 42892 40468 42944 40477
rect 46664 40505 46716 40520
rect 46664 40471 46709 40505
rect 46709 40471 46716 40505
rect 46664 40468 46716 40471
rect 42708 40400 42760 40452
rect 45192 40400 45244 40452
rect 46480 40443 46532 40452
rect 46480 40409 46489 40443
rect 46489 40409 46523 40443
rect 46523 40409 46532 40443
rect 46480 40400 46532 40409
rect 46572 40443 46624 40452
rect 46572 40409 46581 40443
rect 46581 40409 46615 40443
rect 46615 40409 46624 40443
rect 47584 40604 47636 40656
rect 47860 40604 47912 40656
rect 47400 40511 47452 40520
rect 47400 40477 47409 40511
rect 47409 40477 47443 40511
rect 47443 40477 47452 40511
rect 47400 40468 47452 40477
rect 48412 40536 48464 40588
rect 47860 40511 47912 40520
rect 47860 40477 47869 40511
rect 47869 40477 47903 40511
rect 47903 40477 47912 40511
rect 47860 40468 47912 40477
rect 47952 40468 48004 40520
rect 49332 40468 49384 40520
rect 49884 40604 49936 40656
rect 51540 40604 51592 40656
rect 50068 40536 50120 40588
rect 50528 40536 50580 40588
rect 51632 40579 51684 40588
rect 51632 40545 51641 40579
rect 51641 40545 51675 40579
rect 51675 40545 51684 40579
rect 51632 40536 51684 40545
rect 51448 40468 51500 40520
rect 52736 40468 52788 40520
rect 55496 40511 55548 40520
rect 55496 40477 55505 40511
rect 55505 40477 55539 40511
rect 55539 40477 55548 40511
rect 55496 40468 55548 40477
rect 55772 40511 55824 40520
rect 55772 40477 55781 40511
rect 55781 40477 55815 40511
rect 55815 40477 55824 40511
rect 55772 40468 55824 40477
rect 56416 40468 56468 40520
rect 47492 40443 47544 40452
rect 46572 40400 46624 40409
rect 40408 40332 40460 40384
rect 40592 40332 40644 40384
rect 41512 40332 41564 40384
rect 47492 40409 47501 40443
rect 47501 40409 47535 40443
rect 47535 40409 47544 40443
rect 47492 40400 47544 40409
rect 47676 40443 47728 40452
rect 47676 40409 47711 40443
rect 47711 40409 47728 40443
rect 47676 40400 47728 40409
rect 48136 40400 48188 40452
rect 51172 40400 51224 40452
rect 51264 40332 51316 40384
rect 52184 40400 52236 40452
rect 54760 40400 54812 40452
rect 56232 40400 56284 40452
rect 51908 40375 51960 40384
rect 51908 40341 51917 40375
rect 51917 40341 51951 40375
rect 51951 40341 51960 40375
rect 51908 40332 51960 40341
rect 52460 40332 52512 40384
rect 55312 40375 55364 40384
rect 55312 40341 55321 40375
rect 55321 40341 55355 40375
rect 55355 40341 55364 40375
rect 55312 40332 55364 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 23940 40171 23992 40180
rect 23940 40137 23949 40171
rect 23949 40137 23983 40171
rect 23983 40137 23992 40171
rect 23940 40128 23992 40137
rect 20536 40060 20588 40112
rect 22284 40103 22336 40112
rect 22284 40069 22293 40103
rect 22293 40069 22327 40103
rect 22327 40069 22336 40103
rect 22284 40060 22336 40069
rect 25412 40128 25464 40180
rect 25504 40128 25556 40180
rect 30196 40128 30248 40180
rect 30380 40128 30432 40180
rect 31668 40128 31720 40180
rect 37924 40171 37976 40180
rect 37924 40137 37933 40171
rect 37933 40137 37967 40171
rect 37967 40137 37976 40171
rect 37924 40128 37976 40137
rect 38476 40171 38528 40180
rect 38476 40137 38485 40171
rect 38485 40137 38519 40171
rect 38519 40137 38528 40171
rect 38476 40128 38528 40137
rect 40684 40128 40736 40180
rect 46940 40128 46992 40180
rect 47676 40128 47728 40180
rect 22192 39992 22244 40044
rect 22836 39992 22888 40044
rect 24308 40060 24360 40112
rect 24492 39992 24544 40044
rect 26240 40035 26292 40044
rect 26240 40001 26249 40035
rect 26249 40001 26283 40035
rect 26283 40001 26292 40035
rect 26240 39992 26292 40001
rect 27620 39992 27672 40044
rect 29368 40060 29420 40112
rect 31300 40060 31352 40112
rect 30380 39992 30432 40044
rect 30840 40035 30892 40044
rect 30840 40001 30849 40035
rect 30849 40001 30883 40035
rect 30883 40001 30892 40035
rect 30840 39992 30892 40001
rect 32128 39992 32180 40044
rect 32312 39992 32364 40044
rect 32772 39992 32824 40044
rect 33048 40035 33100 40044
rect 33048 40001 33055 40035
rect 33055 40001 33100 40035
rect 33048 39992 33100 40001
rect 34520 40060 34572 40112
rect 39488 40103 39540 40112
rect 39488 40069 39497 40103
rect 39497 40069 39531 40103
rect 39531 40069 39540 40103
rect 39488 40060 39540 40069
rect 35440 39992 35492 40044
rect 38384 40035 38436 40044
rect 38384 40001 38393 40035
rect 38393 40001 38427 40035
rect 38427 40001 38436 40035
rect 38384 39992 38436 40001
rect 40316 40060 40368 40112
rect 40592 40103 40644 40112
rect 40592 40069 40601 40103
rect 40601 40069 40635 40103
rect 40635 40069 40644 40103
rect 40592 40060 40644 40069
rect 23664 39967 23716 39976
rect 23664 39933 23673 39967
rect 23673 39933 23707 39967
rect 23707 39933 23716 39967
rect 23664 39924 23716 39933
rect 2228 39788 2280 39840
rect 25412 39924 25464 39976
rect 33140 39924 33192 39976
rect 33232 39924 33284 39976
rect 34888 39967 34940 39976
rect 34888 39933 34897 39967
rect 34897 39933 34931 39967
rect 34931 39933 34940 39967
rect 34888 39924 34940 39933
rect 34980 39967 35032 39976
rect 34980 39933 34989 39967
rect 34989 39933 35023 39967
rect 35023 39933 35032 39967
rect 34980 39924 35032 39933
rect 36820 39924 36872 39976
rect 41512 40035 41564 40044
rect 41512 40001 41521 40035
rect 41521 40001 41555 40035
rect 41555 40001 41564 40035
rect 41512 39992 41564 40001
rect 45560 40060 45612 40112
rect 45836 40060 45888 40112
rect 46664 40060 46716 40112
rect 47124 40060 47176 40112
rect 42248 39992 42300 40044
rect 42708 39992 42760 40044
rect 44824 39992 44876 40044
rect 39488 39924 39540 39976
rect 39856 39924 39908 39976
rect 46572 39992 46624 40044
rect 48872 40128 48924 40180
rect 48780 40060 48832 40112
rect 49240 40103 49292 40112
rect 49240 40069 49249 40103
rect 49249 40069 49283 40103
rect 49283 40069 49292 40103
rect 49240 40060 49292 40069
rect 45560 39924 45612 39976
rect 49884 40035 49936 40044
rect 49884 40001 49893 40035
rect 49893 40001 49927 40035
rect 49927 40001 49936 40035
rect 51080 40128 51132 40180
rect 52736 40128 52788 40180
rect 52828 40128 52880 40180
rect 49884 39992 49936 40001
rect 50804 40035 50856 40044
rect 50804 40001 50813 40035
rect 50813 40001 50847 40035
rect 50847 40001 50856 40035
rect 50804 39992 50856 40001
rect 51172 39992 51224 40044
rect 51724 39992 51776 40044
rect 51908 39992 51960 40044
rect 56232 40128 56284 40180
rect 56416 40128 56468 40180
rect 55772 40060 55824 40112
rect 54116 40035 54168 40044
rect 54116 40001 54125 40035
rect 54125 40001 54159 40035
rect 54159 40001 54168 40035
rect 54116 39992 54168 40001
rect 54760 40035 54812 40044
rect 54760 40001 54769 40035
rect 54769 40001 54803 40035
rect 54803 40001 54812 40035
rect 54760 39992 54812 40001
rect 51356 39924 51408 39976
rect 55220 39992 55272 40044
rect 55312 39992 55364 40044
rect 56324 39992 56376 40044
rect 57888 40035 57940 40044
rect 57888 40001 57897 40035
rect 57897 40001 57931 40035
rect 57931 40001 57940 40035
rect 57888 39992 57940 40001
rect 28908 39899 28960 39908
rect 28908 39865 28917 39899
rect 28917 39865 28951 39899
rect 28951 39865 28960 39899
rect 28908 39856 28960 39865
rect 30288 39856 30340 39908
rect 48320 39856 48372 39908
rect 27528 39788 27580 39840
rect 29000 39788 29052 39840
rect 31852 39788 31904 39840
rect 32588 39788 32640 39840
rect 33232 39788 33284 39840
rect 34520 39831 34572 39840
rect 34520 39797 34529 39831
rect 34529 39797 34563 39831
rect 34563 39797 34572 39831
rect 34520 39788 34572 39797
rect 40132 39788 40184 39840
rect 41420 39788 41472 39840
rect 44180 39788 44232 39840
rect 44364 39788 44416 39840
rect 45100 39788 45152 39840
rect 45376 39831 45428 39840
rect 45376 39797 45385 39831
rect 45385 39797 45419 39831
rect 45419 39797 45428 39831
rect 45376 39788 45428 39797
rect 45560 39788 45612 39840
rect 46480 39788 46532 39840
rect 47492 39788 47544 39840
rect 49332 39831 49384 39840
rect 49332 39797 49341 39831
rect 49341 39797 49375 39831
rect 49375 39797 49384 39831
rect 49332 39788 49384 39797
rect 55128 39967 55180 39976
rect 55128 39933 55137 39967
rect 55137 39933 55171 39967
rect 55171 39933 55180 39967
rect 55128 39924 55180 39933
rect 56416 39924 56468 39976
rect 52828 39856 52880 39908
rect 53932 39856 53984 39908
rect 53196 39831 53248 39840
rect 53196 39797 53205 39831
rect 53205 39797 53239 39831
rect 53239 39797 53248 39831
rect 53196 39788 53248 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 24308 39584 24360 39636
rect 24492 39584 24544 39636
rect 24584 39584 24636 39636
rect 33048 39584 33100 39636
rect 23940 39516 23992 39568
rect 3884 39380 3936 39432
rect 4620 39380 4672 39432
rect 20904 39423 20956 39432
rect 20904 39389 20913 39423
rect 20913 39389 20947 39423
rect 20947 39389 20956 39423
rect 20904 39380 20956 39389
rect 21916 39448 21968 39500
rect 24124 39448 24176 39500
rect 22744 39423 22796 39432
rect 22744 39389 22753 39423
rect 22753 39389 22787 39423
rect 22787 39389 22796 39423
rect 22744 39380 22796 39389
rect 24584 39380 24636 39432
rect 29828 39516 29880 39568
rect 32128 39516 32180 39568
rect 33692 39516 33744 39568
rect 28908 39448 28960 39500
rect 24860 39423 24912 39432
rect 24860 39389 24874 39423
rect 24874 39389 24908 39423
rect 24908 39389 24912 39423
rect 24860 39380 24912 39389
rect 25044 39423 25096 39432
rect 25044 39389 25053 39423
rect 25053 39389 25087 39423
rect 25087 39389 25096 39423
rect 25044 39380 25096 39389
rect 25504 39380 25556 39432
rect 27528 39380 27580 39432
rect 27896 39423 27948 39432
rect 27896 39389 27930 39423
rect 27930 39389 27948 39423
rect 27896 39380 27948 39389
rect 30196 39380 30248 39432
rect 31484 39380 31536 39432
rect 31760 39423 31812 39432
rect 31760 39389 31769 39423
rect 31769 39389 31803 39423
rect 31803 39389 31812 39423
rect 31760 39380 31812 39389
rect 32128 39423 32180 39432
rect 23848 39312 23900 39364
rect 2412 39244 2464 39296
rect 21088 39287 21140 39296
rect 21088 39253 21097 39287
rect 21097 39253 21131 39287
rect 21131 39253 21140 39287
rect 21088 39244 21140 39253
rect 27620 39244 27672 39296
rect 30288 39244 30340 39296
rect 32128 39389 32137 39423
rect 32137 39389 32171 39423
rect 32171 39389 32180 39423
rect 32128 39380 32180 39389
rect 32496 39380 32548 39432
rect 32588 39312 32640 39364
rect 32220 39244 32272 39296
rect 32404 39287 32456 39296
rect 32404 39253 32413 39287
rect 32413 39253 32447 39287
rect 32447 39253 32456 39287
rect 32404 39244 32456 39253
rect 32772 39380 32824 39432
rect 33140 39423 33192 39432
rect 33140 39389 33149 39423
rect 33149 39389 33183 39423
rect 33183 39389 33192 39423
rect 33140 39380 33192 39389
rect 33324 39423 33376 39432
rect 33324 39389 33357 39423
rect 33357 39389 33376 39423
rect 33324 39380 33376 39389
rect 34336 39312 34388 39364
rect 34796 39448 34848 39500
rect 34888 39423 34940 39432
rect 34888 39389 34897 39423
rect 34897 39389 34931 39423
rect 34931 39389 34940 39423
rect 34888 39380 34940 39389
rect 39580 39584 39632 39636
rect 40132 39584 40184 39636
rect 40960 39584 41012 39636
rect 41604 39584 41656 39636
rect 41880 39584 41932 39636
rect 44364 39584 44416 39636
rect 35440 39516 35492 39568
rect 45192 39584 45244 39636
rect 45284 39584 45336 39636
rect 47216 39584 47268 39636
rect 54116 39584 54168 39636
rect 55496 39584 55548 39636
rect 56416 39627 56468 39636
rect 56416 39593 56425 39627
rect 56425 39593 56459 39627
rect 56459 39593 56468 39627
rect 56416 39584 56468 39593
rect 56784 39627 56836 39636
rect 56784 39593 56793 39627
rect 56793 39593 56827 39627
rect 56827 39593 56836 39627
rect 56784 39584 56836 39593
rect 45008 39516 45060 39568
rect 45560 39516 45612 39568
rect 46664 39516 46716 39568
rect 49332 39516 49384 39568
rect 55220 39516 55272 39568
rect 38660 39448 38712 39500
rect 40408 39448 40460 39500
rect 37280 39380 37332 39432
rect 39304 39380 39356 39432
rect 40040 39380 40092 39432
rect 40224 39380 40276 39432
rect 45008 39380 45060 39432
rect 45284 39423 45336 39432
rect 45284 39389 45293 39423
rect 45293 39389 45327 39423
rect 45327 39389 45336 39423
rect 45284 39380 45336 39389
rect 45652 39423 45704 39432
rect 33324 39244 33376 39296
rect 33508 39287 33560 39296
rect 33508 39253 33517 39287
rect 33517 39253 33551 39287
rect 33551 39253 33560 39287
rect 33508 39244 33560 39253
rect 34612 39244 34664 39296
rect 35808 39312 35860 39364
rect 39948 39312 40000 39364
rect 40592 39312 40644 39364
rect 40868 39355 40920 39364
rect 40868 39321 40877 39355
rect 40877 39321 40911 39355
rect 40911 39321 40920 39355
rect 44088 39355 44140 39364
rect 40868 39312 40920 39321
rect 44088 39321 44097 39355
rect 44097 39321 44131 39355
rect 44131 39321 44140 39355
rect 44088 39312 44140 39321
rect 44824 39312 44876 39364
rect 45192 39312 45244 39364
rect 45652 39389 45661 39423
rect 45661 39389 45695 39423
rect 45695 39389 45704 39423
rect 45652 39380 45704 39389
rect 35992 39244 36044 39296
rect 37372 39244 37424 39296
rect 37740 39244 37792 39296
rect 38568 39244 38620 39296
rect 44732 39244 44784 39296
rect 45100 39244 45152 39296
rect 51172 39491 51224 39500
rect 51172 39457 51181 39491
rect 51181 39457 51215 39491
rect 51215 39457 51224 39491
rect 51172 39448 51224 39457
rect 54484 39491 54536 39500
rect 54484 39457 54493 39491
rect 54493 39457 54527 39491
rect 54527 39457 54536 39491
rect 54484 39448 54536 39457
rect 48596 39423 48648 39432
rect 48596 39389 48605 39423
rect 48605 39389 48639 39423
rect 48639 39389 48648 39423
rect 48596 39380 48648 39389
rect 48688 39423 48740 39432
rect 48688 39389 48697 39423
rect 48697 39389 48731 39423
rect 48731 39389 48740 39423
rect 48964 39423 49016 39432
rect 48688 39380 48740 39389
rect 48964 39389 48973 39423
rect 48973 39389 49007 39423
rect 49007 39389 49016 39423
rect 48964 39380 49016 39389
rect 51632 39380 51684 39432
rect 53656 39380 53708 39432
rect 56324 39423 56376 39432
rect 56324 39389 56333 39423
rect 56333 39389 56367 39423
rect 56367 39389 56376 39423
rect 56324 39380 56376 39389
rect 57796 39380 57848 39432
rect 50068 39312 50120 39364
rect 47216 39244 47268 39296
rect 49424 39244 49476 39296
rect 50804 39244 50856 39296
rect 51172 39244 51224 39296
rect 57336 39287 57388 39296
rect 57336 39253 57345 39287
rect 57345 39253 57379 39287
rect 57379 39253 57388 39287
rect 57336 39244 57388 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 23388 39040 23440 39092
rect 28908 39040 28960 39092
rect 29092 39040 29144 39092
rect 29828 39040 29880 39092
rect 2412 39015 2464 39024
rect 2412 38981 2421 39015
rect 2421 38981 2455 39015
rect 2455 38981 2464 39015
rect 2412 38972 2464 38981
rect 22836 38972 22888 39024
rect 2228 38947 2280 38956
rect 2228 38913 2237 38947
rect 2237 38913 2271 38947
rect 2271 38913 2280 38947
rect 2228 38904 2280 38913
rect 2780 38879 2832 38888
rect 2780 38845 2789 38879
rect 2789 38845 2823 38879
rect 2823 38845 2832 38879
rect 2780 38836 2832 38845
rect 21088 38947 21140 38956
rect 21088 38913 21097 38947
rect 21097 38913 21131 38947
rect 21131 38913 21140 38947
rect 21088 38904 21140 38913
rect 21180 38836 21232 38888
rect 22100 38904 22152 38956
rect 22376 38904 22428 38956
rect 22652 38904 22704 38956
rect 22284 38879 22336 38888
rect 22284 38845 22293 38879
rect 22293 38845 22327 38879
rect 22327 38845 22336 38879
rect 23388 38904 23440 38956
rect 23848 38947 23900 38956
rect 23848 38913 23857 38947
rect 23857 38913 23891 38947
rect 23891 38913 23900 38947
rect 23848 38904 23900 38913
rect 27620 38904 27672 38956
rect 29552 38904 29604 38956
rect 30012 38904 30064 38956
rect 30196 38904 30248 38956
rect 22284 38836 22336 38845
rect 20996 38768 21048 38820
rect 23204 38768 23256 38820
rect 24400 38836 24452 38888
rect 24676 38836 24728 38888
rect 23848 38768 23900 38820
rect 30472 38972 30524 39024
rect 30748 39083 30800 39092
rect 30748 39049 30773 39083
rect 30773 39049 30800 39083
rect 30748 39040 30800 39049
rect 31024 39040 31076 39092
rect 31484 39083 31536 39092
rect 31484 39049 31493 39083
rect 31493 39049 31527 39083
rect 31527 39049 31536 39083
rect 31484 39040 31536 39049
rect 33048 39083 33100 39092
rect 33048 39049 33057 39083
rect 33057 39049 33091 39083
rect 33091 39049 33100 39083
rect 33048 39040 33100 39049
rect 35440 39040 35492 39092
rect 30840 38904 30892 38956
rect 31760 38972 31812 39024
rect 32312 38972 32364 39024
rect 32680 39015 32732 39024
rect 32680 38981 32689 39015
rect 32689 38981 32723 39015
rect 32723 38981 32732 39015
rect 32680 38972 32732 38981
rect 36084 38972 36136 39024
rect 32496 38947 32548 38956
rect 32496 38913 32506 38947
rect 32506 38913 32540 38947
rect 32540 38913 32548 38947
rect 32496 38904 32548 38913
rect 33324 38904 33376 38956
rect 33784 38904 33836 38956
rect 34888 38904 34940 38956
rect 37280 38947 37332 38956
rect 34152 38836 34204 38888
rect 32496 38768 32548 38820
rect 33600 38811 33652 38820
rect 33600 38777 33609 38811
rect 33609 38777 33643 38811
rect 33643 38777 33652 38811
rect 33600 38768 33652 38777
rect 34244 38768 34296 38820
rect 19524 38700 19576 38752
rect 20812 38700 20864 38752
rect 22192 38743 22244 38752
rect 22192 38709 22201 38743
rect 22201 38709 22235 38743
rect 22235 38709 22244 38743
rect 22192 38700 22244 38709
rect 22928 38743 22980 38752
rect 22928 38709 22937 38743
rect 22937 38709 22971 38743
rect 22971 38709 22980 38743
rect 23940 38743 23992 38752
rect 22928 38700 22980 38709
rect 23940 38709 23949 38743
rect 23949 38709 23983 38743
rect 23983 38709 23992 38743
rect 23940 38700 23992 38709
rect 30012 38700 30064 38752
rect 30932 38743 30984 38752
rect 30932 38709 30941 38743
rect 30941 38709 30975 38743
rect 30975 38709 30984 38743
rect 30932 38700 30984 38709
rect 35716 38836 35768 38888
rect 37280 38913 37289 38947
rect 37289 38913 37323 38947
rect 37323 38913 37332 38947
rect 37280 38904 37332 38913
rect 37648 39040 37700 39092
rect 38476 39040 38528 39092
rect 40224 39040 40276 39092
rect 40500 39040 40552 39092
rect 45652 39040 45704 39092
rect 46020 39040 46072 39092
rect 49240 39040 49292 39092
rect 52092 39083 52144 39092
rect 52092 39049 52101 39083
rect 52101 39049 52135 39083
rect 52135 39049 52144 39083
rect 52092 39040 52144 39049
rect 53472 39083 53524 39092
rect 53472 39049 53481 39083
rect 53481 39049 53515 39083
rect 53515 39049 53524 39083
rect 53472 39040 53524 39049
rect 39396 38972 39448 39024
rect 37832 38904 37884 38956
rect 38384 38947 38436 38956
rect 38384 38913 38393 38947
rect 38393 38913 38427 38947
rect 38427 38913 38436 38947
rect 38384 38904 38436 38913
rect 38568 38947 38620 38956
rect 38568 38913 38577 38947
rect 38577 38913 38611 38947
rect 38611 38913 38620 38947
rect 38568 38904 38620 38913
rect 39488 38836 39540 38888
rect 40040 38947 40092 38956
rect 40040 38913 40049 38947
rect 40049 38913 40083 38947
rect 40083 38913 40092 38947
rect 40040 38904 40092 38913
rect 41604 38972 41656 39024
rect 42156 38972 42208 39024
rect 40592 38947 40644 38956
rect 40592 38913 40601 38947
rect 40601 38913 40635 38947
rect 40635 38913 40644 38947
rect 40592 38904 40644 38913
rect 41512 38947 41564 38956
rect 41512 38913 41521 38947
rect 41521 38913 41555 38947
rect 41555 38913 41564 38947
rect 41512 38904 41564 38913
rect 35624 38768 35676 38820
rect 39028 38768 39080 38820
rect 39396 38768 39448 38820
rect 39672 38768 39724 38820
rect 40132 38768 40184 38820
rect 43536 38836 43588 38888
rect 34336 38700 34388 38752
rect 34796 38700 34848 38752
rect 35532 38700 35584 38752
rect 37648 38700 37700 38752
rect 40592 38743 40644 38752
rect 40592 38709 40601 38743
rect 40601 38709 40635 38743
rect 40635 38709 40644 38743
rect 40592 38700 40644 38709
rect 45376 38972 45428 39024
rect 44364 38904 44416 38956
rect 44732 38947 44784 38956
rect 44732 38913 44741 38947
rect 44741 38913 44775 38947
rect 44775 38913 44784 38947
rect 44732 38904 44784 38913
rect 45008 38947 45060 38956
rect 45008 38913 45017 38947
rect 45017 38913 45051 38947
rect 45051 38913 45060 38947
rect 45008 38904 45060 38913
rect 44088 38836 44140 38888
rect 45468 38904 45520 38956
rect 45836 38904 45888 38956
rect 48504 39015 48556 39024
rect 48504 38981 48513 39015
rect 48513 38981 48547 39015
rect 48547 38981 48556 39015
rect 48504 38972 48556 38981
rect 48780 38972 48832 39024
rect 45560 38836 45612 38888
rect 48044 38904 48096 38956
rect 44732 38768 44784 38820
rect 46296 38768 46348 38820
rect 44272 38700 44324 38752
rect 44456 38743 44508 38752
rect 44456 38709 44465 38743
rect 44465 38709 44499 38743
rect 44499 38709 44508 38743
rect 44456 38700 44508 38709
rect 44640 38700 44692 38752
rect 45744 38700 45796 38752
rect 46940 38836 46992 38888
rect 48412 38836 48464 38888
rect 48964 38836 49016 38888
rect 49700 38836 49752 38888
rect 49884 38836 49936 38888
rect 50620 38904 50672 38956
rect 50712 38879 50764 38888
rect 50712 38845 50721 38879
rect 50721 38845 50755 38879
rect 50755 38845 50764 38879
rect 50712 38836 50764 38845
rect 52184 38947 52236 38956
rect 51908 38836 51960 38888
rect 46940 38743 46992 38752
rect 46940 38709 46949 38743
rect 46949 38709 46983 38743
rect 46983 38709 46992 38743
rect 46940 38700 46992 38709
rect 48688 38700 48740 38752
rect 48964 38700 49016 38752
rect 52184 38913 52193 38947
rect 52193 38913 52227 38947
rect 52227 38913 52236 38947
rect 52184 38904 52236 38913
rect 53288 38947 53340 38956
rect 53288 38913 53297 38947
rect 53297 38913 53331 38947
rect 53331 38913 53340 38947
rect 53288 38904 53340 38913
rect 53656 38836 53708 38888
rect 51448 38700 51500 38752
rect 51724 38700 51776 38752
rect 56600 38700 56652 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 21180 38496 21232 38548
rect 20628 38292 20680 38344
rect 19524 38267 19576 38276
rect 19524 38233 19558 38267
rect 19558 38233 19576 38267
rect 19524 38224 19576 38233
rect 23940 38496 23992 38548
rect 29368 38496 29420 38548
rect 22284 38428 22336 38480
rect 24400 38428 24452 38480
rect 26700 38471 26752 38480
rect 24584 38360 24636 38412
rect 26700 38437 26709 38471
rect 26709 38437 26743 38471
rect 26743 38437 26752 38471
rect 26700 38428 26752 38437
rect 27528 38428 27580 38480
rect 27712 38428 27764 38480
rect 30288 38428 30340 38480
rect 34796 38496 34848 38548
rect 36728 38496 36780 38548
rect 22376 38292 22428 38344
rect 22652 38292 22704 38344
rect 22928 38335 22980 38344
rect 22928 38301 22937 38335
rect 22937 38301 22971 38335
rect 22971 38301 22980 38335
rect 22928 38292 22980 38301
rect 23204 38335 23256 38344
rect 23204 38301 23213 38335
rect 23213 38301 23247 38335
rect 23247 38301 23256 38335
rect 23204 38292 23256 38301
rect 24492 38292 24544 38344
rect 25044 38335 25096 38344
rect 25044 38301 25053 38335
rect 25053 38301 25087 38335
rect 25087 38301 25096 38335
rect 25044 38292 25096 38301
rect 28540 38292 28592 38344
rect 30932 38360 30984 38412
rect 31116 38360 31168 38412
rect 22468 38224 22520 38276
rect 26516 38267 26568 38276
rect 26516 38233 26525 38267
rect 26525 38233 26559 38267
rect 26559 38233 26568 38267
rect 26516 38224 26568 38233
rect 30380 38292 30432 38344
rect 30472 38292 30524 38344
rect 30748 38292 30800 38344
rect 30104 38224 30156 38276
rect 20720 38156 20772 38208
rect 21640 38199 21692 38208
rect 21640 38165 21649 38199
rect 21649 38165 21683 38199
rect 21683 38165 21692 38199
rect 21640 38156 21692 38165
rect 22100 38156 22152 38208
rect 22652 38156 22704 38208
rect 25504 38156 25556 38208
rect 29828 38156 29880 38208
rect 31484 38224 31536 38276
rect 33324 38292 33376 38344
rect 34152 38292 34204 38344
rect 35164 38403 35216 38412
rect 35164 38369 35173 38403
rect 35173 38369 35207 38403
rect 35207 38369 35216 38403
rect 35164 38360 35216 38369
rect 31300 38156 31352 38208
rect 34336 38156 34388 38208
rect 34612 38156 34664 38208
rect 34796 38156 34848 38208
rect 35624 38292 35676 38344
rect 36268 38292 36320 38344
rect 36544 38360 36596 38412
rect 37556 38428 37608 38480
rect 38660 38496 38712 38548
rect 41328 38496 41380 38548
rect 44732 38496 44784 38548
rect 46112 38496 46164 38548
rect 46296 38539 46348 38548
rect 46296 38505 46305 38539
rect 46305 38505 46339 38539
rect 46339 38505 46348 38539
rect 46296 38496 46348 38505
rect 49976 38496 50028 38548
rect 51632 38539 51684 38548
rect 51632 38505 51641 38539
rect 51641 38505 51675 38539
rect 51675 38505 51684 38539
rect 51632 38496 51684 38505
rect 52184 38496 52236 38548
rect 38752 38403 38804 38412
rect 36636 38335 36688 38344
rect 36636 38301 36645 38335
rect 36645 38301 36679 38335
rect 36679 38301 36688 38335
rect 38752 38369 38761 38403
rect 38761 38369 38795 38403
rect 38795 38369 38804 38403
rect 38752 38360 38804 38369
rect 39672 38428 39724 38480
rect 41696 38428 41748 38480
rect 44364 38428 44416 38480
rect 46204 38428 46256 38480
rect 46388 38428 46440 38480
rect 49056 38428 49108 38480
rect 53288 38496 53340 38548
rect 53656 38539 53708 38548
rect 53656 38505 53665 38539
rect 53665 38505 53699 38539
rect 53699 38505 53708 38539
rect 53656 38496 53708 38505
rect 40040 38360 40092 38412
rect 42432 38360 42484 38412
rect 45192 38360 45244 38412
rect 36636 38292 36688 38301
rect 37280 38292 37332 38344
rect 37832 38335 37884 38344
rect 37832 38301 37841 38335
rect 37841 38301 37875 38335
rect 37875 38301 37884 38335
rect 37832 38292 37884 38301
rect 39856 38335 39908 38344
rect 36728 38267 36780 38276
rect 36728 38233 36737 38267
rect 36737 38233 36771 38267
rect 36771 38233 36780 38267
rect 36728 38224 36780 38233
rect 37556 38224 37608 38276
rect 38476 38224 38528 38276
rect 35900 38156 35952 38208
rect 37096 38156 37148 38208
rect 39856 38301 39865 38335
rect 39865 38301 39899 38335
rect 39899 38301 39908 38335
rect 39856 38292 39908 38301
rect 39948 38292 40000 38344
rect 40684 38335 40736 38344
rect 40684 38301 40693 38335
rect 40693 38301 40727 38335
rect 40727 38301 40736 38335
rect 40684 38292 40736 38301
rect 41512 38335 41564 38344
rect 39028 38224 39080 38276
rect 41512 38301 41521 38335
rect 41521 38301 41555 38335
rect 41555 38301 41564 38335
rect 41512 38292 41564 38301
rect 41604 38224 41656 38276
rect 38936 38156 38988 38208
rect 40316 38156 40368 38208
rect 41236 38156 41288 38208
rect 44456 38292 44508 38344
rect 46020 38292 46072 38344
rect 46388 38292 46440 38344
rect 43536 38267 43588 38276
rect 43536 38233 43545 38267
rect 43545 38233 43579 38267
rect 43579 38233 43588 38267
rect 43536 38224 43588 38233
rect 43720 38267 43772 38276
rect 43720 38233 43755 38267
rect 43755 38233 43772 38267
rect 43720 38224 43772 38233
rect 46296 38224 46348 38276
rect 46664 38295 46670 38322
rect 46670 38295 46704 38322
rect 46704 38295 46716 38322
rect 46664 38270 46716 38295
rect 46756 38335 46808 38344
rect 46756 38301 46770 38335
rect 46770 38301 46804 38335
rect 46804 38301 46808 38335
rect 46756 38292 46808 38301
rect 46940 38335 46992 38344
rect 46940 38301 46949 38335
rect 46949 38301 46983 38335
rect 46983 38301 46992 38335
rect 46940 38292 46992 38301
rect 48412 38292 48464 38344
rect 48872 38292 48924 38344
rect 51080 38360 51132 38412
rect 53748 38403 53800 38412
rect 47492 38267 47544 38276
rect 47492 38233 47501 38267
rect 47501 38233 47535 38267
rect 47535 38233 47544 38267
rect 47492 38224 47544 38233
rect 49700 38292 49752 38344
rect 53748 38369 53757 38403
rect 53757 38369 53791 38403
rect 53791 38369 53800 38403
rect 53748 38360 53800 38369
rect 56600 38360 56652 38412
rect 57888 38403 57940 38412
rect 57888 38369 57897 38403
rect 57897 38369 57931 38403
rect 57931 38369 57940 38403
rect 57888 38360 57940 38369
rect 53012 38292 53064 38344
rect 50712 38224 50764 38276
rect 51448 38267 51500 38276
rect 51448 38233 51457 38267
rect 51457 38233 51491 38267
rect 51491 38233 51500 38267
rect 51448 38224 51500 38233
rect 51540 38224 51592 38276
rect 57336 38224 57388 38276
rect 44824 38156 44876 38208
rect 46204 38156 46256 38208
rect 48320 38156 48372 38208
rect 56784 38156 56836 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 22468 37952 22520 38004
rect 22652 37995 22704 38004
rect 22652 37961 22661 37995
rect 22661 37961 22695 37995
rect 22695 37961 22704 37995
rect 22652 37952 22704 37961
rect 24584 37995 24636 38004
rect 24584 37961 24593 37995
rect 24593 37961 24627 37995
rect 24627 37961 24636 37995
rect 24584 37952 24636 37961
rect 24676 37995 24728 38004
rect 24676 37961 24685 37995
rect 24685 37961 24719 37995
rect 24719 37961 24728 37995
rect 24676 37952 24728 37961
rect 20720 37816 20772 37868
rect 20536 37748 20588 37800
rect 22376 37791 22428 37800
rect 22376 37757 22385 37791
rect 22385 37757 22419 37791
rect 22419 37757 22428 37791
rect 22376 37748 22428 37757
rect 22652 37748 22704 37800
rect 22928 37748 22980 37800
rect 26976 37952 27028 38004
rect 28172 37952 28224 38004
rect 29552 37952 29604 38004
rect 30472 37952 30524 38004
rect 31116 37952 31168 38004
rect 32588 37952 32640 38004
rect 32956 37952 33008 38004
rect 30196 37884 30248 37936
rect 24492 37859 24544 37868
rect 24492 37825 24501 37859
rect 24501 37825 24535 37859
rect 24535 37825 24544 37859
rect 24492 37816 24544 37825
rect 25044 37816 25096 37868
rect 20352 37612 20404 37664
rect 20996 37612 21048 37664
rect 22836 37612 22888 37664
rect 25504 37655 25556 37664
rect 25504 37621 25513 37655
rect 25513 37621 25547 37655
rect 25547 37621 25556 37655
rect 25504 37612 25556 37621
rect 30748 37859 30800 37868
rect 30748 37825 30757 37859
rect 30757 37825 30791 37859
rect 30791 37825 30800 37859
rect 30748 37816 30800 37825
rect 34152 37816 34204 37868
rect 30012 37791 30064 37800
rect 26240 37680 26292 37732
rect 30012 37757 30021 37791
rect 30021 37757 30055 37791
rect 30055 37757 30064 37791
rect 30012 37748 30064 37757
rect 30104 37791 30156 37800
rect 30104 37757 30113 37791
rect 30113 37757 30147 37791
rect 30147 37757 30156 37791
rect 31024 37791 31076 37800
rect 30104 37748 30156 37757
rect 31024 37757 31033 37791
rect 31033 37757 31067 37791
rect 31067 37757 31076 37791
rect 31024 37748 31076 37757
rect 32588 37791 32640 37800
rect 31300 37680 31352 37732
rect 32588 37757 32597 37791
rect 32597 37757 32631 37791
rect 32631 37757 32640 37791
rect 32588 37748 32640 37757
rect 33140 37748 33192 37800
rect 33324 37748 33376 37800
rect 35808 37884 35860 37936
rect 35716 37816 35768 37868
rect 33784 37680 33836 37732
rect 26148 37655 26200 37664
rect 26148 37621 26157 37655
rect 26157 37621 26191 37655
rect 26191 37621 26200 37655
rect 26148 37612 26200 37621
rect 34060 37612 34112 37664
rect 34152 37612 34204 37664
rect 36268 37952 36320 38004
rect 39580 37952 39632 38004
rect 39948 37995 40000 38004
rect 39948 37961 39957 37995
rect 39957 37961 39991 37995
rect 39991 37961 40000 37995
rect 39948 37952 40000 37961
rect 41236 37995 41288 38004
rect 41236 37961 41245 37995
rect 41245 37961 41279 37995
rect 41279 37961 41288 37995
rect 41236 37952 41288 37961
rect 36636 37884 36688 37936
rect 36176 37859 36228 37868
rect 36176 37825 36205 37859
rect 36205 37825 36228 37859
rect 36452 37859 36504 37868
rect 36176 37816 36228 37825
rect 36452 37825 36461 37859
rect 36461 37825 36495 37859
rect 36495 37825 36504 37859
rect 36452 37816 36504 37825
rect 37832 37884 37884 37936
rect 39488 37884 39540 37936
rect 39764 37884 39816 37936
rect 40684 37884 40736 37936
rect 41144 37884 41196 37936
rect 43536 37952 43588 38004
rect 45376 37952 45428 38004
rect 46756 37952 46808 38004
rect 47124 37952 47176 38004
rect 49700 37952 49752 38004
rect 52184 37995 52236 38004
rect 52184 37961 52193 37995
rect 52193 37961 52227 37995
rect 52227 37961 52236 37995
rect 52184 37952 52236 37961
rect 40132 37859 40184 37868
rect 37188 37748 37240 37800
rect 37372 37748 37424 37800
rect 37556 37680 37608 37732
rect 40132 37825 40141 37859
rect 40141 37825 40175 37859
rect 40175 37825 40184 37859
rect 40132 37816 40184 37825
rect 40316 37816 40368 37868
rect 40408 37816 40460 37868
rect 50712 37884 50764 37936
rect 51908 37884 51960 37936
rect 41604 37816 41656 37868
rect 42064 37816 42116 37868
rect 42432 37859 42484 37868
rect 42432 37825 42441 37859
rect 42441 37825 42475 37859
rect 42475 37825 42484 37859
rect 42432 37816 42484 37825
rect 42800 37816 42852 37868
rect 43536 37816 43588 37868
rect 42156 37748 42208 37800
rect 45560 37816 45612 37868
rect 46112 37816 46164 37868
rect 46480 37859 46532 37868
rect 46480 37825 46489 37859
rect 46489 37825 46523 37859
rect 46523 37825 46532 37859
rect 46480 37816 46532 37825
rect 47216 37816 47268 37868
rect 47676 37816 47728 37868
rect 48596 37816 48648 37868
rect 44732 37748 44784 37800
rect 45836 37748 45888 37800
rect 46204 37748 46256 37800
rect 46388 37748 46440 37800
rect 49056 37816 49108 37868
rect 49516 37816 49568 37868
rect 49792 37859 49844 37868
rect 49792 37825 49801 37859
rect 49801 37825 49835 37859
rect 49835 37825 49844 37859
rect 49792 37816 49844 37825
rect 49976 37859 50028 37868
rect 49976 37825 49985 37859
rect 49985 37825 50019 37859
rect 50019 37825 50028 37859
rect 49976 37816 50028 37825
rect 50068 37859 50120 37868
rect 50068 37825 50077 37859
rect 50077 37825 50111 37859
rect 50111 37825 50120 37859
rect 50068 37816 50120 37825
rect 50252 37816 50304 37868
rect 50620 37816 50672 37868
rect 52184 37816 52236 37868
rect 56784 37859 56836 37868
rect 56784 37825 56793 37859
rect 56793 37825 56827 37859
rect 56827 37825 56836 37859
rect 56784 37816 56836 37825
rect 49884 37748 49936 37800
rect 53196 37791 53248 37800
rect 45652 37680 45704 37732
rect 47400 37680 47452 37732
rect 48872 37680 48924 37732
rect 50620 37680 50672 37732
rect 36728 37655 36780 37664
rect 36728 37621 36737 37655
rect 36737 37621 36771 37655
rect 36771 37621 36780 37655
rect 36728 37612 36780 37621
rect 37464 37612 37516 37664
rect 41052 37612 41104 37664
rect 47860 37612 47912 37664
rect 48136 37612 48188 37664
rect 50160 37612 50212 37664
rect 53196 37757 53205 37791
rect 53205 37757 53239 37791
rect 53239 37757 53248 37791
rect 53196 37748 53248 37757
rect 56876 37791 56928 37800
rect 56876 37757 56885 37791
rect 56885 37757 56919 37791
rect 56919 37757 56928 37791
rect 56876 37748 56928 37757
rect 57152 37791 57204 37800
rect 57152 37757 57161 37791
rect 57161 37757 57195 37791
rect 57195 37757 57204 37791
rect 57152 37748 57204 37757
rect 53932 37680 53984 37732
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 20904 37408 20956 37460
rect 23388 37451 23440 37460
rect 23388 37417 23397 37451
rect 23397 37417 23431 37451
rect 23431 37417 23440 37451
rect 23388 37408 23440 37417
rect 26516 37408 26568 37460
rect 27252 37408 27304 37460
rect 30380 37408 30432 37460
rect 31116 37408 31168 37460
rect 20812 37272 20864 37324
rect 31300 37272 31352 37324
rect 32312 37272 32364 37324
rect 34152 37408 34204 37460
rect 34336 37408 34388 37460
rect 33784 37340 33836 37392
rect 33416 37272 33468 37324
rect 36452 37408 36504 37460
rect 39304 37408 39356 37460
rect 37372 37340 37424 37392
rect 20352 37247 20404 37256
rect 20352 37213 20361 37247
rect 20361 37213 20395 37247
rect 20395 37213 20404 37247
rect 20352 37204 20404 37213
rect 20628 37204 20680 37256
rect 21640 37179 21692 37188
rect 21640 37145 21674 37179
rect 21674 37145 21692 37179
rect 21640 37136 21692 37145
rect 22376 37204 22428 37256
rect 26700 37204 26752 37256
rect 29644 37204 29696 37256
rect 30012 37204 30064 37256
rect 31024 37204 31076 37256
rect 31208 37204 31260 37256
rect 31484 37204 31536 37256
rect 31852 37204 31904 37256
rect 34796 37272 34848 37324
rect 36360 37272 36412 37324
rect 26148 37179 26200 37188
rect 26148 37145 26182 37179
rect 26182 37145 26200 37179
rect 26148 37136 26200 37145
rect 30288 37179 30340 37188
rect 30288 37145 30297 37179
rect 30297 37145 30331 37179
rect 30331 37145 30340 37179
rect 30288 37136 30340 37145
rect 31668 37136 31720 37188
rect 35716 37204 35768 37256
rect 36084 37204 36136 37256
rect 22376 37068 22428 37120
rect 26240 37068 26292 37120
rect 31852 37068 31904 37120
rect 32128 37111 32180 37120
rect 32128 37077 32137 37111
rect 32137 37077 32171 37111
rect 32171 37077 32180 37111
rect 32128 37068 32180 37077
rect 33968 37136 34020 37188
rect 37556 37272 37608 37324
rect 37280 37204 37332 37256
rect 38752 37340 38804 37392
rect 40592 37408 40644 37460
rect 42064 37408 42116 37460
rect 42156 37408 42208 37460
rect 44732 37408 44784 37460
rect 45192 37408 45244 37460
rect 46020 37408 46072 37460
rect 47400 37451 47452 37460
rect 41420 37340 41472 37392
rect 42708 37340 42760 37392
rect 46388 37340 46440 37392
rect 47400 37417 47409 37451
rect 47409 37417 47443 37451
rect 47443 37417 47452 37451
rect 47400 37408 47452 37417
rect 47860 37451 47912 37460
rect 47860 37417 47869 37451
rect 47869 37417 47903 37451
rect 47903 37417 47912 37451
rect 47860 37408 47912 37417
rect 48136 37340 48188 37392
rect 56048 37340 56100 37392
rect 40408 37204 40460 37256
rect 40592 37247 40644 37256
rect 40592 37213 40601 37247
rect 40601 37213 40635 37247
rect 40635 37213 40644 37247
rect 40592 37204 40644 37213
rect 44732 37272 44784 37324
rect 41052 37204 41104 37256
rect 41144 37204 41196 37256
rect 42432 37204 42484 37256
rect 45376 37272 45428 37324
rect 46296 37272 46348 37324
rect 47216 37272 47268 37324
rect 49056 37272 49108 37324
rect 45284 37204 45336 37256
rect 46112 37247 46164 37256
rect 34796 37068 34848 37120
rect 36176 37068 36228 37120
rect 38384 37111 38436 37120
rect 38384 37077 38393 37111
rect 38393 37077 38427 37111
rect 38427 37077 38436 37111
rect 38384 37068 38436 37077
rect 40592 37068 40644 37120
rect 42156 37136 42208 37188
rect 46112 37213 46121 37247
rect 46121 37213 46155 37247
rect 46155 37213 46164 37247
rect 46112 37204 46164 37213
rect 46204 37247 46256 37256
rect 46204 37213 46213 37247
rect 46213 37213 46247 37247
rect 46247 37213 46256 37247
rect 46204 37204 46256 37213
rect 46480 37204 46532 37256
rect 47492 37204 47544 37256
rect 48136 37247 48188 37256
rect 48136 37213 48145 37247
rect 48145 37213 48179 37247
rect 48179 37213 48188 37247
rect 48136 37204 48188 37213
rect 48504 37204 48556 37256
rect 49516 37272 49568 37324
rect 49700 37272 49752 37324
rect 51264 37272 51316 37324
rect 51816 37272 51868 37324
rect 56600 37315 56652 37324
rect 56600 37281 56609 37315
rect 56609 37281 56643 37315
rect 56643 37281 56652 37315
rect 56600 37272 56652 37281
rect 50252 37204 50304 37256
rect 41512 37068 41564 37120
rect 43444 37111 43496 37120
rect 43444 37077 43453 37111
rect 43453 37077 43487 37111
rect 43487 37077 43496 37111
rect 43444 37068 43496 37077
rect 44456 37068 44508 37120
rect 45652 37068 45704 37120
rect 48320 37136 48372 37188
rect 48412 37136 48464 37188
rect 50620 37247 50672 37256
rect 50620 37213 50629 37247
rect 50629 37213 50663 37247
rect 50663 37213 50672 37247
rect 50620 37204 50672 37213
rect 57980 37204 58032 37256
rect 47676 37068 47728 37120
rect 48136 37068 48188 37120
rect 57152 37136 57204 37188
rect 49976 37068 50028 37120
rect 52184 37068 52236 37120
rect 56784 37068 56836 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 24492 36864 24544 36916
rect 22560 36796 22612 36848
rect 31668 36864 31720 36916
rect 31852 36864 31904 36916
rect 32220 36864 32272 36916
rect 32956 36864 33008 36916
rect 33140 36864 33192 36916
rect 44824 36907 44876 36916
rect 22376 36728 22428 36780
rect 22836 36771 22888 36780
rect 22836 36737 22845 36771
rect 22845 36737 22879 36771
rect 22879 36737 22888 36771
rect 22836 36728 22888 36737
rect 22928 36771 22980 36780
rect 22928 36737 22937 36771
rect 22937 36737 22971 36771
rect 22971 36737 22980 36771
rect 22928 36728 22980 36737
rect 22192 36660 22244 36712
rect 26332 36660 26384 36712
rect 29368 36771 29420 36780
rect 29368 36737 29377 36771
rect 29377 36737 29411 36771
rect 29411 36737 29420 36771
rect 29368 36728 29420 36737
rect 29644 36796 29696 36848
rect 32404 36728 32456 36780
rect 33416 36771 33468 36780
rect 33416 36737 33425 36771
rect 33425 36737 33459 36771
rect 33459 36737 33468 36771
rect 33416 36728 33468 36737
rect 34152 36796 34204 36848
rect 33784 36728 33836 36780
rect 23204 36592 23256 36644
rect 28632 36660 28684 36712
rect 29000 36660 29052 36712
rect 29276 36660 29328 36712
rect 34336 36703 34388 36712
rect 34336 36669 34345 36703
rect 34345 36669 34379 36703
rect 34379 36669 34388 36703
rect 34336 36660 34388 36669
rect 34796 36660 34848 36712
rect 35808 36796 35860 36848
rect 36360 36839 36412 36848
rect 36360 36805 36369 36839
rect 36369 36805 36403 36839
rect 36403 36805 36412 36839
rect 36360 36796 36412 36805
rect 37740 36796 37792 36848
rect 40408 36796 40460 36848
rect 40592 36796 40644 36848
rect 41144 36796 41196 36848
rect 41420 36796 41472 36848
rect 35256 36771 35308 36780
rect 35256 36737 35265 36771
rect 35265 36737 35299 36771
rect 35299 36737 35308 36771
rect 35256 36728 35308 36737
rect 35624 36728 35676 36780
rect 36176 36771 36228 36780
rect 36176 36737 36185 36771
rect 36185 36737 36219 36771
rect 36219 36737 36228 36771
rect 36176 36728 36228 36737
rect 36452 36771 36504 36780
rect 36452 36737 36461 36771
rect 36461 36737 36495 36771
rect 36495 36737 36504 36771
rect 36452 36728 36504 36737
rect 36544 36771 36596 36780
rect 36544 36737 36553 36771
rect 36553 36737 36587 36771
rect 36587 36737 36596 36771
rect 36544 36728 36596 36737
rect 25136 36524 25188 36576
rect 26608 36524 26660 36576
rect 27804 36524 27856 36576
rect 29828 36524 29880 36576
rect 30472 36524 30524 36576
rect 30656 36524 30708 36576
rect 32864 36592 32916 36644
rect 33968 36592 34020 36644
rect 35256 36592 35308 36644
rect 35716 36660 35768 36712
rect 37372 36728 37424 36780
rect 40500 36728 40552 36780
rect 44456 36771 44508 36780
rect 44456 36737 44465 36771
rect 44465 36737 44499 36771
rect 44499 36737 44508 36771
rect 44456 36728 44508 36737
rect 35992 36592 36044 36644
rect 42708 36592 42760 36644
rect 44824 36873 44833 36907
rect 44833 36873 44867 36907
rect 44867 36873 44876 36907
rect 44824 36864 44876 36873
rect 48596 36839 48648 36848
rect 48596 36805 48605 36839
rect 48605 36805 48639 36839
rect 48639 36805 48648 36839
rect 48596 36796 48648 36805
rect 49148 36796 49200 36848
rect 49792 36839 49844 36848
rect 49792 36805 49801 36839
rect 49801 36805 49835 36839
rect 49835 36805 49844 36839
rect 49792 36796 49844 36805
rect 45836 36728 45888 36780
rect 46756 36728 46808 36780
rect 48780 36728 48832 36780
rect 50068 36796 50120 36848
rect 56600 36864 56652 36916
rect 56876 36864 56928 36916
rect 57980 36907 58032 36916
rect 50160 36728 50212 36780
rect 54024 36771 54076 36780
rect 54024 36737 54033 36771
rect 54033 36737 54067 36771
rect 54067 36737 54076 36771
rect 54024 36728 54076 36737
rect 47492 36660 47544 36712
rect 48136 36660 48188 36712
rect 49608 36660 49660 36712
rect 53932 36703 53984 36712
rect 53932 36669 53941 36703
rect 53941 36669 53975 36703
rect 53975 36669 53984 36703
rect 53932 36660 53984 36669
rect 46940 36592 46992 36644
rect 56508 36728 56560 36780
rect 57244 36728 57296 36780
rect 57980 36873 57989 36907
rect 57989 36873 58023 36907
rect 58023 36873 58032 36907
rect 57980 36864 58032 36873
rect 54944 36703 54996 36712
rect 54944 36669 54953 36703
rect 54953 36669 54987 36703
rect 54987 36669 54996 36703
rect 54944 36660 54996 36669
rect 57336 36592 57388 36644
rect 57612 36592 57664 36644
rect 33508 36524 33560 36576
rect 34796 36524 34848 36576
rect 35624 36524 35676 36576
rect 37372 36524 37424 36576
rect 37832 36567 37884 36576
rect 37832 36533 37841 36567
rect 37841 36533 37875 36567
rect 37875 36533 37884 36567
rect 37832 36524 37884 36533
rect 44640 36567 44692 36576
rect 44640 36533 44649 36567
rect 44649 36533 44683 36567
rect 44683 36533 44692 36567
rect 44640 36524 44692 36533
rect 48044 36524 48096 36576
rect 48964 36524 49016 36576
rect 49424 36524 49476 36576
rect 49976 36567 50028 36576
rect 49976 36533 49985 36567
rect 49985 36533 50019 36567
rect 50019 36533 50028 36567
rect 49976 36524 50028 36533
rect 52276 36524 52328 36576
rect 57152 36567 57204 36576
rect 57152 36533 57161 36567
rect 57161 36533 57195 36567
rect 57195 36533 57204 36567
rect 57152 36524 57204 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 26608 36363 26660 36372
rect 26608 36329 26617 36363
rect 26617 36329 26651 36363
rect 26651 36329 26660 36363
rect 26608 36320 26660 36329
rect 31576 36320 31628 36372
rect 34152 36320 34204 36372
rect 34520 36320 34572 36372
rect 35716 36363 35768 36372
rect 33876 36252 33928 36304
rect 29828 36227 29880 36236
rect 29828 36193 29837 36227
rect 29837 36193 29871 36227
rect 29871 36193 29880 36227
rect 29828 36184 29880 36193
rect 25044 36116 25096 36168
rect 26056 36048 26108 36100
rect 26700 36159 26752 36168
rect 26700 36125 26709 36159
rect 26709 36125 26743 36159
rect 26743 36125 26752 36159
rect 27528 36159 27580 36168
rect 26700 36116 26752 36125
rect 27528 36125 27537 36159
rect 27537 36125 27571 36159
rect 27571 36125 27580 36159
rect 27528 36116 27580 36125
rect 27804 36159 27856 36168
rect 27804 36125 27838 36159
rect 27838 36125 27856 36159
rect 27804 36116 27856 36125
rect 31024 36116 31076 36168
rect 34704 36184 34756 36236
rect 34980 36252 35032 36304
rect 35716 36329 35725 36363
rect 35725 36329 35759 36363
rect 35759 36329 35768 36363
rect 35716 36320 35768 36329
rect 36452 36320 36504 36372
rect 40316 36320 40368 36372
rect 43444 36363 43496 36372
rect 43444 36329 43453 36363
rect 43453 36329 43487 36363
rect 43487 36329 43496 36363
rect 43444 36320 43496 36329
rect 45560 36363 45612 36372
rect 45560 36329 45569 36363
rect 45569 36329 45603 36363
rect 45603 36329 45612 36363
rect 45560 36320 45612 36329
rect 54944 36320 54996 36372
rect 56416 36363 56468 36372
rect 56416 36329 56425 36363
rect 56425 36329 56459 36363
rect 56459 36329 56468 36363
rect 56416 36320 56468 36329
rect 57244 36363 57296 36372
rect 57244 36329 57253 36363
rect 57253 36329 57287 36363
rect 57287 36329 57296 36363
rect 57244 36320 57296 36329
rect 32864 36159 32916 36168
rect 32864 36125 32873 36159
rect 32873 36125 32907 36159
rect 32907 36125 32916 36159
rect 32864 36116 32916 36125
rect 33968 36159 34020 36168
rect 33968 36125 33977 36159
rect 33977 36125 34011 36159
rect 34011 36125 34020 36159
rect 33968 36116 34020 36125
rect 25504 35980 25556 36032
rect 26240 36023 26292 36032
rect 26240 35989 26249 36023
rect 26249 35989 26283 36023
rect 26283 35989 26292 36023
rect 26240 35980 26292 35989
rect 28632 35980 28684 36032
rect 32128 36048 32180 36100
rect 33232 36048 33284 36100
rect 34520 36116 34572 36168
rect 34796 36116 34848 36168
rect 37280 36252 37332 36304
rect 35256 36116 35308 36168
rect 36084 36184 36136 36236
rect 48044 36227 48096 36236
rect 36820 36116 36872 36168
rect 43168 36159 43220 36168
rect 43168 36125 43177 36159
rect 43177 36125 43211 36159
rect 43211 36125 43220 36159
rect 43168 36116 43220 36125
rect 44272 36159 44324 36168
rect 44272 36125 44281 36159
rect 44281 36125 44315 36159
rect 44315 36125 44324 36159
rect 44272 36116 44324 36125
rect 45284 36116 45336 36168
rect 46112 36159 46164 36168
rect 46112 36125 46121 36159
rect 46121 36125 46155 36159
rect 46155 36125 46164 36159
rect 46112 36116 46164 36125
rect 46204 36116 46256 36168
rect 48044 36193 48053 36227
rect 48053 36193 48087 36227
rect 48087 36193 48096 36227
rect 48044 36184 48096 36193
rect 52276 36227 52328 36236
rect 52276 36193 52285 36227
rect 52285 36193 52319 36227
rect 52319 36193 52328 36227
rect 52276 36184 52328 36193
rect 56140 36227 56192 36236
rect 56140 36193 56149 36227
rect 56149 36193 56183 36227
rect 56183 36193 56192 36227
rect 56140 36184 56192 36193
rect 57060 36184 57112 36236
rect 48228 36159 48280 36168
rect 48228 36125 48237 36159
rect 48237 36125 48271 36159
rect 48271 36125 48280 36159
rect 48228 36116 48280 36125
rect 52368 36159 52420 36168
rect 32404 35980 32456 36032
rect 34796 35980 34848 36032
rect 35992 36048 36044 36100
rect 45468 36048 45520 36100
rect 46940 36048 46992 36100
rect 47676 36048 47728 36100
rect 52368 36125 52377 36159
rect 52377 36125 52411 36159
rect 52411 36125 52420 36159
rect 52368 36116 52420 36125
rect 56048 36159 56100 36168
rect 52092 36048 52144 36100
rect 56048 36125 56057 36159
rect 56057 36125 56091 36159
rect 56091 36125 56100 36159
rect 56048 36116 56100 36125
rect 56968 36048 57020 36100
rect 41696 35980 41748 36032
rect 43536 35980 43588 36032
rect 44456 35980 44508 36032
rect 47492 35980 47544 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 26056 35776 26108 35828
rect 26240 35708 26292 35760
rect 25044 35683 25096 35692
rect 25044 35649 25053 35683
rect 25053 35649 25087 35683
rect 25087 35649 25096 35683
rect 25044 35640 25096 35649
rect 25596 35640 25648 35692
rect 30380 35708 30432 35760
rect 30748 35708 30800 35760
rect 30932 35708 30984 35760
rect 31944 35708 31996 35760
rect 32864 35708 32916 35760
rect 34980 35708 35032 35760
rect 35808 35776 35860 35828
rect 43168 35776 43220 35828
rect 43904 35776 43956 35828
rect 44364 35776 44416 35828
rect 46204 35776 46256 35828
rect 48596 35776 48648 35828
rect 26608 35504 26660 35556
rect 26700 35436 26752 35488
rect 29000 35640 29052 35692
rect 31852 35640 31904 35692
rect 33968 35640 34020 35692
rect 35256 35640 35308 35692
rect 38752 35708 38804 35760
rect 37372 35640 37424 35692
rect 40408 35683 40460 35692
rect 40408 35649 40417 35683
rect 40417 35649 40451 35683
rect 40451 35649 40460 35683
rect 40408 35640 40460 35649
rect 43352 35708 43404 35760
rect 43444 35751 43496 35760
rect 43444 35717 43453 35751
rect 43453 35717 43487 35751
rect 43487 35717 43496 35751
rect 43444 35708 43496 35717
rect 31484 35615 31536 35624
rect 31484 35581 31493 35615
rect 31493 35581 31527 35615
rect 31527 35581 31536 35615
rect 31484 35572 31536 35581
rect 32956 35572 33008 35624
rect 33048 35504 33100 35556
rect 35532 35572 35584 35624
rect 37280 35615 37332 35624
rect 37280 35581 37289 35615
rect 37289 35581 37323 35615
rect 37323 35581 37332 35615
rect 37280 35572 37332 35581
rect 41512 35572 41564 35624
rect 41696 35615 41748 35624
rect 41696 35581 41705 35615
rect 41705 35581 41739 35615
rect 41739 35581 41748 35615
rect 41696 35572 41748 35581
rect 43536 35640 43588 35692
rect 45192 35708 45244 35760
rect 46296 35708 46348 35760
rect 49332 35708 49384 35760
rect 49884 35708 49936 35760
rect 51172 35708 51224 35760
rect 56784 35708 56836 35760
rect 44088 35640 44140 35692
rect 44272 35683 44324 35692
rect 44272 35649 44281 35683
rect 44281 35649 44315 35683
rect 44315 35649 44324 35683
rect 44272 35640 44324 35649
rect 44456 35683 44508 35692
rect 44456 35649 44465 35683
rect 44465 35649 44499 35683
rect 44499 35649 44508 35683
rect 44456 35640 44508 35649
rect 45008 35640 45060 35692
rect 46388 35640 46440 35692
rect 48412 35640 48464 35692
rect 49240 35640 49292 35692
rect 50712 35683 50764 35692
rect 50712 35649 50721 35683
rect 50721 35649 50755 35683
rect 50755 35649 50764 35683
rect 50712 35640 50764 35649
rect 51448 35683 51500 35692
rect 51448 35649 51457 35683
rect 51457 35649 51491 35683
rect 51491 35649 51500 35683
rect 51448 35640 51500 35649
rect 56140 35683 56192 35692
rect 44364 35572 44416 35624
rect 46112 35572 46164 35624
rect 48596 35572 48648 35624
rect 51632 35572 51684 35624
rect 36176 35504 36228 35556
rect 56140 35649 56149 35683
rect 56149 35649 56183 35683
rect 56183 35649 56192 35683
rect 56140 35640 56192 35649
rect 29276 35479 29328 35488
rect 29276 35445 29285 35479
rect 29285 35445 29319 35479
rect 29319 35445 29328 35479
rect 29276 35436 29328 35445
rect 33232 35436 33284 35488
rect 34152 35479 34204 35488
rect 34152 35445 34161 35479
rect 34161 35445 34195 35479
rect 34195 35445 34204 35479
rect 34152 35436 34204 35445
rect 35992 35436 36044 35488
rect 38752 35436 38804 35488
rect 40960 35436 41012 35488
rect 41328 35436 41380 35488
rect 42892 35479 42944 35488
rect 42892 35445 42901 35479
rect 42901 35445 42935 35479
rect 42935 35445 42944 35479
rect 42892 35436 42944 35445
rect 43628 35436 43680 35488
rect 45100 35479 45152 35488
rect 45100 35445 45109 35479
rect 45109 35445 45143 35479
rect 45143 35445 45152 35479
rect 45100 35436 45152 35445
rect 49056 35436 49108 35488
rect 50160 35479 50212 35488
rect 50160 35445 50169 35479
rect 50169 35445 50203 35479
rect 50203 35445 50212 35479
rect 50160 35436 50212 35445
rect 50620 35436 50672 35488
rect 53380 35436 53432 35488
rect 56048 35436 56100 35488
rect 56324 35436 56376 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 25044 35232 25096 35284
rect 27528 35232 27580 35284
rect 30012 35232 30064 35284
rect 32588 35232 32640 35284
rect 41052 35232 41104 35284
rect 41880 35275 41932 35284
rect 41880 35241 41889 35275
rect 41889 35241 41923 35275
rect 41923 35241 41932 35275
rect 41880 35232 41932 35241
rect 42708 35232 42760 35284
rect 47216 35275 47268 35284
rect 26332 35164 26384 35216
rect 30932 35164 30984 35216
rect 28172 35139 28224 35148
rect 28172 35105 28181 35139
rect 28181 35105 28215 35139
rect 28215 35105 28224 35139
rect 28172 35096 28224 35105
rect 30748 35096 30800 35148
rect 31024 35139 31076 35148
rect 31024 35105 31033 35139
rect 31033 35105 31067 35139
rect 31067 35105 31076 35139
rect 31024 35096 31076 35105
rect 34704 35139 34756 35148
rect 34704 35105 34713 35139
rect 34713 35105 34747 35139
rect 34747 35105 34756 35139
rect 34704 35096 34756 35105
rect 40960 35139 41012 35148
rect 40960 35105 40969 35139
rect 40969 35105 41003 35139
rect 41003 35105 41012 35139
rect 40960 35096 41012 35105
rect 41052 35139 41104 35148
rect 41052 35105 41061 35139
rect 41061 35105 41095 35139
rect 41095 35105 41104 35139
rect 41052 35096 41104 35105
rect 42524 35096 42576 35148
rect 25136 35071 25188 35080
rect 25136 35037 25170 35071
rect 25170 35037 25188 35071
rect 25136 35028 25188 35037
rect 27252 35071 27304 35080
rect 27252 35037 27261 35071
rect 27261 35037 27295 35071
rect 27295 35037 27304 35071
rect 27252 35028 27304 35037
rect 27620 35028 27672 35080
rect 30840 35028 30892 35080
rect 37280 35028 37332 35080
rect 37832 35028 37884 35080
rect 38660 35028 38712 35080
rect 31944 34960 31996 35012
rect 35440 34960 35492 35012
rect 41328 35028 41380 35080
rect 42892 35164 42944 35216
rect 43352 35096 43404 35148
rect 43628 35139 43680 35148
rect 43628 35105 43637 35139
rect 43637 35105 43671 35139
rect 43671 35105 43680 35139
rect 43628 35096 43680 35105
rect 45100 35096 45152 35148
rect 45468 35164 45520 35216
rect 47216 35241 47225 35275
rect 47225 35241 47259 35275
rect 47259 35241 47268 35275
rect 47216 35232 47268 35241
rect 49056 35232 49108 35284
rect 52092 35232 52144 35284
rect 52368 35232 52420 35284
rect 57152 35232 57204 35284
rect 48688 35164 48740 35216
rect 51172 35164 51224 35216
rect 52276 35164 52328 35216
rect 51264 35139 51316 35148
rect 51264 35105 51273 35139
rect 51273 35105 51307 35139
rect 51307 35105 51316 35139
rect 51264 35096 51316 35105
rect 52552 35139 52604 35148
rect 52552 35105 52561 35139
rect 52561 35105 52595 35139
rect 52595 35105 52604 35139
rect 52552 35096 52604 35105
rect 44272 35028 44324 35080
rect 45008 35028 45060 35080
rect 30104 34892 30156 34944
rect 37188 34892 37240 34944
rect 39120 34892 39172 34944
rect 43260 34960 43312 35012
rect 43720 34960 43772 35012
rect 44916 34960 44968 35012
rect 41420 34892 41472 34944
rect 45928 34960 45980 35012
rect 46388 35071 46440 35080
rect 46388 35037 46397 35071
rect 46397 35037 46431 35071
rect 46431 35037 46440 35071
rect 46388 35028 46440 35037
rect 47216 35028 47268 35080
rect 46296 34935 46348 34944
rect 46296 34901 46305 34935
rect 46305 34901 46339 34935
rect 46339 34901 46348 34935
rect 46296 34892 46348 34901
rect 47400 34960 47452 35012
rect 48964 34960 49016 35012
rect 49976 35028 50028 35080
rect 50160 35028 50212 35080
rect 52460 35071 52512 35080
rect 52460 35037 52469 35071
rect 52469 35037 52503 35071
rect 52503 35037 52512 35071
rect 52460 35028 52512 35037
rect 52644 35071 52696 35080
rect 52644 35037 52653 35071
rect 52653 35037 52687 35071
rect 52687 35037 52696 35071
rect 52644 35028 52696 35037
rect 53380 35071 53432 35080
rect 53380 35037 53389 35071
rect 53389 35037 53423 35071
rect 53423 35037 53432 35071
rect 53380 35028 53432 35037
rect 56324 35028 56376 35080
rect 56968 35071 57020 35080
rect 51172 34935 51224 34944
rect 51172 34901 51181 34935
rect 51181 34901 51215 34935
rect 51215 34901 51224 34935
rect 51172 34892 51224 34901
rect 52460 34892 52512 34944
rect 52736 34892 52788 34944
rect 55588 34960 55640 35012
rect 56968 35037 56977 35071
rect 56977 35037 57011 35071
rect 57011 35037 57020 35071
rect 56968 35028 57020 35037
rect 57060 35071 57112 35080
rect 57060 35037 57069 35071
rect 57069 35037 57103 35071
rect 57103 35037 57112 35071
rect 57060 35028 57112 35037
rect 53472 34892 53524 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 31852 34688 31904 34740
rect 38660 34731 38712 34740
rect 38660 34697 38669 34731
rect 38669 34697 38703 34731
rect 38703 34697 38712 34731
rect 38660 34688 38712 34697
rect 40408 34688 40460 34740
rect 30380 34620 30432 34672
rect 28172 34595 28224 34604
rect 28172 34561 28181 34595
rect 28181 34561 28215 34595
rect 28215 34561 28224 34595
rect 28172 34552 28224 34561
rect 27620 34484 27672 34536
rect 27712 34348 27764 34400
rect 32312 34595 32364 34604
rect 32312 34561 32321 34595
rect 32321 34561 32355 34595
rect 32355 34561 32364 34595
rect 32588 34595 32640 34604
rect 32312 34552 32364 34561
rect 32588 34561 32597 34595
rect 32597 34561 32631 34595
rect 32631 34561 32640 34595
rect 32588 34552 32640 34561
rect 33232 34595 33284 34604
rect 33232 34561 33241 34595
rect 33241 34561 33275 34595
rect 33275 34561 33284 34595
rect 33232 34552 33284 34561
rect 35716 34620 35768 34672
rect 34152 34552 34204 34604
rect 38384 34620 38436 34672
rect 40316 34620 40368 34672
rect 41328 34620 41380 34672
rect 41512 34688 41564 34740
rect 44364 34731 44416 34740
rect 42800 34620 42852 34672
rect 42892 34620 42944 34672
rect 44364 34697 44373 34731
rect 44373 34697 44407 34731
rect 44407 34697 44416 34731
rect 44364 34688 44416 34697
rect 44456 34688 44508 34740
rect 49884 34688 49936 34740
rect 49976 34688 50028 34740
rect 40408 34595 40460 34604
rect 31484 34484 31536 34536
rect 31944 34416 31996 34468
rect 35532 34484 35584 34536
rect 40408 34561 40417 34595
rect 40417 34561 40451 34595
rect 40451 34561 40460 34595
rect 40408 34552 40460 34561
rect 41420 34552 41472 34604
rect 41512 34595 41564 34604
rect 41512 34561 41521 34595
rect 41521 34561 41555 34595
rect 41555 34561 41564 34595
rect 41512 34552 41564 34561
rect 43352 34552 43404 34604
rect 44180 34595 44232 34604
rect 44180 34561 44189 34595
rect 44189 34561 44223 34595
rect 44223 34561 44232 34595
rect 44180 34552 44232 34561
rect 44456 34552 44508 34604
rect 45100 34552 45152 34604
rect 45192 34595 45244 34604
rect 45192 34561 45201 34595
rect 45201 34561 45235 34595
rect 45235 34561 45244 34595
rect 47492 34620 47544 34672
rect 45192 34552 45244 34561
rect 40500 34484 40552 34536
rect 43352 34416 43404 34468
rect 44824 34484 44876 34536
rect 45468 34484 45520 34536
rect 45192 34416 45244 34468
rect 47124 34552 47176 34604
rect 46940 34527 46992 34536
rect 46940 34493 46949 34527
rect 46949 34493 46983 34527
rect 46983 34493 46992 34527
rect 46940 34484 46992 34493
rect 47676 34552 47728 34604
rect 48412 34552 48464 34604
rect 48688 34552 48740 34604
rect 49056 34595 49108 34604
rect 49056 34561 49065 34595
rect 49065 34561 49099 34595
rect 49099 34561 49108 34595
rect 49056 34552 49108 34561
rect 47308 34484 47360 34536
rect 49240 34484 49292 34536
rect 50252 34620 50304 34672
rect 50988 34688 51040 34740
rect 51724 34688 51776 34740
rect 52276 34688 52328 34740
rect 50804 34663 50856 34672
rect 50804 34629 50813 34663
rect 50813 34629 50847 34663
rect 50847 34629 50856 34663
rect 50804 34620 50856 34629
rect 49884 34595 49936 34604
rect 49884 34561 49893 34595
rect 49893 34561 49927 34595
rect 49927 34561 49936 34595
rect 49884 34552 49936 34561
rect 50160 34552 50212 34604
rect 51172 34552 51224 34604
rect 51448 34552 51500 34604
rect 51724 34595 51776 34604
rect 51724 34561 51733 34595
rect 51733 34561 51767 34595
rect 51767 34561 51776 34595
rect 51724 34552 51776 34561
rect 52000 34595 52052 34604
rect 52000 34561 52009 34595
rect 52009 34561 52043 34595
rect 52043 34561 52052 34595
rect 52000 34552 52052 34561
rect 52184 34552 52236 34604
rect 56692 34552 56744 34604
rect 53656 34484 53708 34536
rect 41972 34348 42024 34400
rect 44180 34391 44232 34400
rect 44180 34357 44189 34391
rect 44189 34357 44223 34391
rect 44223 34357 44232 34391
rect 44180 34348 44232 34357
rect 44732 34348 44784 34400
rect 45008 34348 45060 34400
rect 46940 34348 46992 34400
rect 47952 34348 48004 34400
rect 48228 34348 48280 34400
rect 50804 34348 50856 34400
rect 51080 34391 51132 34400
rect 51080 34357 51089 34391
rect 51089 34357 51123 34391
rect 51123 34357 51132 34391
rect 51080 34348 51132 34357
rect 56968 34391 57020 34400
rect 56968 34357 56977 34391
rect 56977 34357 57011 34391
rect 57011 34357 57020 34391
rect 56968 34348 57020 34357
rect 58072 34391 58124 34400
rect 58072 34357 58081 34391
rect 58081 34357 58115 34391
rect 58115 34357 58124 34391
rect 58072 34348 58124 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 28172 34187 28224 34196
rect 28172 34153 28181 34187
rect 28181 34153 28215 34187
rect 28215 34153 28224 34187
rect 28172 34144 28224 34153
rect 39120 34187 39172 34196
rect 39120 34153 39129 34187
rect 39129 34153 39163 34187
rect 39163 34153 39172 34187
rect 39120 34144 39172 34153
rect 40132 34144 40184 34196
rect 43904 34144 43956 34196
rect 45008 34144 45060 34196
rect 46296 34144 46348 34196
rect 47492 34144 47544 34196
rect 47584 34144 47636 34196
rect 25504 34051 25556 34060
rect 25504 34017 25513 34051
rect 25513 34017 25547 34051
rect 25547 34017 25556 34051
rect 25504 34008 25556 34017
rect 28632 34051 28684 34060
rect 28632 34017 28641 34051
rect 28641 34017 28675 34051
rect 28675 34017 28684 34051
rect 28632 34008 28684 34017
rect 27712 33983 27764 33992
rect 27712 33949 27721 33983
rect 27721 33949 27755 33983
rect 27755 33949 27764 33983
rect 27712 33940 27764 33949
rect 26056 33872 26108 33924
rect 26884 33872 26936 33924
rect 30104 34008 30156 34060
rect 30380 34008 30432 34060
rect 34704 34051 34756 34060
rect 34704 34017 34713 34051
rect 34713 34017 34747 34051
rect 34747 34017 34756 34051
rect 34704 34008 34756 34017
rect 38660 34008 38712 34060
rect 41052 34008 41104 34060
rect 41604 34008 41656 34060
rect 41972 34051 42024 34060
rect 41972 34017 41981 34051
rect 41981 34017 42015 34051
rect 42015 34017 42024 34051
rect 41972 34008 42024 34017
rect 43812 34076 43864 34128
rect 44272 34119 44324 34128
rect 44272 34085 44281 34119
rect 44281 34085 44315 34119
rect 44315 34085 44324 34119
rect 44272 34076 44324 34085
rect 44180 34051 44232 34060
rect 44180 34017 44189 34051
rect 44189 34017 44223 34051
rect 44223 34017 44232 34051
rect 44180 34008 44232 34017
rect 34612 33940 34664 33992
rect 38752 33940 38804 33992
rect 39120 33940 39172 33992
rect 41880 33983 41932 33992
rect 41880 33949 41889 33983
rect 41889 33949 41923 33983
rect 41923 33949 41932 33983
rect 41880 33940 41932 33949
rect 42984 33940 43036 33992
rect 44916 33940 44968 33992
rect 45100 33940 45152 33992
rect 45744 34076 45796 34128
rect 46940 34008 46992 34060
rect 47216 34008 47268 34060
rect 48320 34008 48372 34060
rect 46480 33983 46532 33992
rect 46480 33949 46489 33983
rect 46489 33949 46523 33983
rect 46523 33949 46532 33983
rect 46480 33940 46532 33949
rect 47400 33983 47452 33992
rect 47400 33949 47409 33983
rect 47409 33949 47443 33983
rect 47443 33949 47452 33983
rect 47400 33940 47452 33949
rect 30748 33872 30800 33924
rect 42524 33872 42576 33924
rect 45008 33915 45060 33924
rect 45008 33881 45017 33915
rect 45017 33881 45051 33915
rect 45051 33881 45060 33915
rect 45008 33872 45060 33881
rect 45376 33872 45428 33924
rect 47308 33872 47360 33924
rect 24124 33804 24176 33856
rect 27528 33847 27580 33856
rect 27528 33813 27537 33847
rect 27537 33813 27571 33847
rect 27571 33813 27580 33847
rect 27528 33804 27580 33813
rect 29092 33804 29144 33856
rect 29920 33804 29972 33856
rect 36084 33847 36136 33856
rect 36084 33813 36093 33847
rect 36093 33813 36127 33847
rect 36127 33813 36136 33847
rect 36084 33804 36136 33813
rect 39304 33847 39356 33856
rect 39304 33813 39313 33847
rect 39313 33813 39347 33847
rect 39347 33813 39356 33847
rect 39304 33804 39356 33813
rect 40684 33847 40736 33856
rect 40684 33813 40693 33847
rect 40693 33813 40727 33847
rect 40727 33813 40736 33847
rect 40684 33804 40736 33813
rect 40868 33804 40920 33856
rect 41236 33804 41288 33856
rect 42800 33847 42852 33856
rect 42800 33813 42809 33847
rect 42809 33813 42843 33847
rect 42843 33813 42852 33847
rect 42800 33804 42852 33813
rect 46940 33804 46992 33856
rect 47216 33804 47268 33856
rect 47860 33940 47912 33992
rect 48412 33983 48464 33992
rect 48412 33949 48421 33983
rect 48421 33949 48455 33983
rect 48455 33949 48464 33983
rect 48412 33940 48464 33949
rect 48412 33804 48464 33856
rect 51356 34144 51408 34196
rect 51632 34144 51684 34196
rect 52644 34144 52696 34196
rect 54484 34187 54536 34196
rect 54484 34153 54493 34187
rect 54493 34153 54527 34187
rect 54527 34153 54536 34187
rect 54484 34144 54536 34153
rect 56140 34144 56192 34196
rect 51632 34008 51684 34060
rect 52552 34008 52604 34060
rect 52736 34008 52788 34060
rect 53472 34051 53524 34060
rect 49884 33940 49936 33992
rect 50068 33940 50120 33992
rect 49332 33915 49384 33924
rect 49332 33881 49341 33915
rect 49341 33881 49375 33915
rect 49375 33881 49384 33915
rect 49332 33872 49384 33881
rect 50160 33872 50212 33924
rect 50896 33940 50948 33992
rect 52368 33940 52420 33992
rect 52460 33940 52512 33992
rect 53472 34017 53481 34051
rect 53481 34017 53515 34051
rect 53515 34017 53524 34051
rect 53472 34008 53524 34017
rect 58072 34076 58124 34128
rect 56968 34008 57020 34060
rect 57888 34051 57940 34060
rect 57888 34017 57897 34051
rect 57897 34017 57931 34051
rect 57931 34017 57940 34051
rect 57888 34008 57940 34017
rect 54484 33983 54536 33992
rect 52184 33872 52236 33924
rect 54484 33949 54493 33983
rect 54493 33949 54527 33983
rect 54527 33949 54536 33983
rect 54484 33940 54536 33949
rect 54668 33983 54720 33992
rect 54668 33949 54677 33983
rect 54677 33949 54711 33983
rect 54711 33949 54720 33983
rect 54668 33940 54720 33949
rect 55588 33983 55640 33992
rect 55588 33949 55597 33983
rect 55597 33949 55631 33983
rect 55631 33949 55640 33983
rect 55588 33940 55640 33949
rect 55864 33940 55916 33992
rect 51356 33804 51408 33856
rect 51724 33804 51776 33856
rect 55496 33804 55548 33856
rect 56324 33804 56376 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 26332 33600 26384 33652
rect 30748 33643 30800 33652
rect 30748 33609 30757 33643
rect 30757 33609 30791 33643
rect 30791 33609 30800 33643
rect 30748 33600 30800 33609
rect 41604 33643 41656 33652
rect 41604 33609 41613 33643
rect 41613 33609 41647 33643
rect 41647 33609 41656 33643
rect 41604 33600 41656 33609
rect 42800 33600 42852 33652
rect 42984 33643 43036 33652
rect 42984 33609 42993 33643
rect 42993 33609 43027 33643
rect 43027 33609 43036 33643
rect 42984 33600 43036 33609
rect 45192 33600 45244 33652
rect 45560 33643 45612 33652
rect 45560 33609 45569 33643
rect 45569 33609 45603 33643
rect 45603 33609 45612 33643
rect 45560 33600 45612 33609
rect 46480 33600 46532 33652
rect 47216 33600 47268 33652
rect 47308 33600 47360 33652
rect 27528 33532 27580 33584
rect 29920 33575 29972 33584
rect 29920 33541 29929 33575
rect 29929 33541 29963 33575
rect 29963 33541 29972 33575
rect 29920 33532 29972 33541
rect 30104 33575 30156 33584
rect 30104 33541 30113 33575
rect 30113 33541 30147 33575
rect 30147 33541 30156 33575
rect 30104 33532 30156 33541
rect 41328 33532 41380 33584
rect 42892 33532 42944 33584
rect 24124 33507 24176 33516
rect 24124 33473 24133 33507
rect 24133 33473 24167 33507
rect 24167 33473 24176 33507
rect 24124 33464 24176 33473
rect 24032 33396 24084 33448
rect 24860 33464 24912 33516
rect 26240 33464 26292 33516
rect 30932 33507 30984 33516
rect 30932 33473 30941 33507
rect 30941 33473 30975 33507
rect 30975 33473 30984 33507
rect 30932 33464 30984 33473
rect 41880 33464 41932 33516
rect 42432 33507 42484 33516
rect 42432 33473 42441 33507
rect 42441 33473 42475 33507
rect 42475 33473 42484 33507
rect 42432 33464 42484 33473
rect 44364 33532 44416 33584
rect 44916 33507 44968 33516
rect 24952 33328 25004 33380
rect 26884 33396 26936 33448
rect 26976 33396 27028 33448
rect 41236 33396 41288 33448
rect 42708 33396 42760 33448
rect 44916 33473 44925 33507
rect 44925 33473 44959 33507
rect 44959 33473 44968 33507
rect 44916 33464 44968 33473
rect 45100 33532 45152 33584
rect 48412 33600 48464 33652
rect 48596 33600 48648 33652
rect 49976 33532 50028 33584
rect 50620 33600 50672 33652
rect 50896 33532 50948 33584
rect 52000 33600 52052 33652
rect 55588 33600 55640 33652
rect 55864 33643 55916 33652
rect 55864 33609 55873 33643
rect 55873 33609 55907 33643
rect 55907 33609 55916 33643
rect 55864 33600 55916 33609
rect 43904 33396 43956 33448
rect 47032 33464 47084 33516
rect 47308 33464 47360 33516
rect 47492 33464 47544 33516
rect 47952 33507 48004 33516
rect 47952 33473 47961 33507
rect 47961 33473 47995 33507
rect 47995 33473 48004 33507
rect 47952 33464 48004 33473
rect 49056 33507 49108 33516
rect 49056 33473 49065 33507
rect 49065 33473 49099 33507
rect 49099 33473 49108 33507
rect 49056 33464 49108 33473
rect 49240 33507 49292 33516
rect 49240 33473 49249 33507
rect 49249 33473 49283 33507
rect 49283 33473 49292 33507
rect 49240 33464 49292 33473
rect 51080 33464 51132 33516
rect 51356 33507 51408 33516
rect 51356 33473 51365 33507
rect 51365 33473 51399 33507
rect 51399 33473 51408 33507
rect 51356 33464 51408 33473
rect 52368 33532 52420 33584
rect 53932 33575 53984 33584
rect 53932 33541 53941 33575
rect 53941 33541 53975 33575
rect 53975 33541 53984 33575
rect 53932 33532 53984 33541
rect 54208 33532 54260 33584
rect 56324 33575 56376 33584
rect 54760 33507 54812 33516
rect 54760 33473 54769 33507
rect 54769 33473 54803 33507
rect 54803 33473 54812 33507
rect 54760 33464 54812 33473
rect 26332 33328 26384 33380
rect 47124 33396 47176 33448
rect 50804 33439 50856 33448
rect 50804 33405 50813 33439
rect 50813 33405 50847 33439
rect 50847 33405 50856 33439
rect 50804 33396 50856 33405
rect 50988 33396 51040 33448
rect 55404 33464 55456 33516
rect 56324 33541 56333 33575
rect 56333 33541 56367 33575
rect 56367 33541 56376 33575
rect 56324 33532 56376 33541
rect 56416 33464 56468 33516
rect 56600 33507 56652 33516
rect 56600 33473 56609 33507
rect 56609 33473 56643 33507
rect 56643 33473 56652 33507
rect 56600 33464 56652 33473
rect 56876 33464 56928 33516
rect 49332 33328 49384 33380
rect 51080 33328 51132 33380
rect 54668 33328 54720 33380
rect 23848 33260 23900 33312
rect 27160 33260 27212 33312
rect 29092 33260 29144 33312
rect 39120 33260 39172 33312
rect 43904 33260 43956 33312
rect 44180 33260 44232 33312
rect 44640 33260 44692 33312
rect 45560 33260 45612 33312
rect 47584 33260 47636 33312
rect 54116 33303 54168 33312
rect 54116 33269 54125 33303
rect 54125 33269 54159 33303
rect 54159 33269 54168 33303
rect 54116 33260 54168 33269
rect 56968 33260 57020 33312
rect 57152 33303 57204 33312
rect 57152 33269 57161 33303
rect 57161 33269 57195 33303
rect 57195 33269 57204 33303
rect 57152 33260 57204 33269
rect 57244 33260 57296 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 26332 33056 26384 33108
rect 41328 33099 41380 33108
rect 41328 33065 41337 33099
rect 41337 33065 41371 33099
rect 41371 33065 41380 33099
rect 41328 33056 41380 33065
rect 42708 33099 42760 33108
rect 42708 33065 42717 33099
rect 42717 33065 42751 33099
rect 42751 33065 42760 33099
rect 42708 33056 42760 33065
rect 44088 33099 44140 33108
rect 44088 33065 44097 33099
rect 44097 33065 44131 33099
rect 44131 33065 44140 33099
rect 44088 33056 44140 33065
rect 44180 33056 44232 33108
rect 44916 33056 44968 33108
rect 45376 33056 45428 33108
rect 46480 33056 46532 33108
rect 46756 33056 46808 33108
rect 47124 33099 47176 33108
rect 47124 33065 47133 33099
rect 47133 33065 47167 33099
rect 47167 33065 47176 33099
rect 47124 33056 47176 33065
rect 29920 32988 29972 33040
rect 26700 32963 26752 32972
rect 26700 32929 26709 32963
rect 26709 32929 26743 32963
rect 26743 32929 26752 32963
rect 26700 32920 26752 32929
rect 26884 32963 26936 32972
rect 26884 32929 26893 32963
rect 26893 32929 26927 32963
rect 26927 32929 26936 32963
rect 26884 32920 26936 32929
rect 26976 32920 27028 32972
rect 30012 32963 30064 32972
rect 30012 32929 30021 32963
rect 30021 32929 30055 32963
rect 30055 32929 30064 32963
rect 30012 32920 30064 32929
rect 30288 32920 30340 32972
rect 23848 32895 23900 32904
rect 23848 32861 23857 32895
rect 23857 32861 23891 32895
rect 23891 32861 23900 32895
rect 23848 32852 23900 32861
rect 25044 32852 25096 32904
rect 35808 32852 35860 32904
rect 37096 32895 37148 32904
rect 37096 32861 37130 32895
rect 37130 32861 37148 32895
rect 37096 32852 37148 32861
rect 41512 32895 41564 32904
rect 41512 32861 41521 32895
rect 41521 32861 41555 32895
rect 41555 32861 41564 32895
rect 41512 32852 41564 32861
rect 41604 32895 41656 32904
rect 41604 32861 41613 32895
rect 41613 32861 41647 32895
rect 41647 32861 41656 32895
rect 42524 32988 42576 33040
rect 48044 33056 48096 33108
rect 48136 33056 48188 33108
rect 50160 33056 50212 33108
rect 51356 33056 51408 33108
rect 54484 33056 54536 33108
rect 55588 33056 55640 33108
rect 56416 33056 56468 33108
rect 44456 32920 44508 32972
rect 41604 32852 41656 32861
rect 28540 32784 28592 32836
rect 41236 32784 41288 32836
rect 44824 32852 44876 32904
rect 45284 32852 45336 32904
rect 47952 32988 48004 33040
rect 51264 33031 51316 33040
rect 51264 32997 51273 33031
rect 51273 32997 51307 33031
rect 51307 32997 51316 33031
rect 51264 32988 51316 32997
rect 46388 32852 46440 32904
rect 26056 32716 26108 32768
rect 27988 32716 28040 32768
rect 29000 32759 29052 32768
rect 29000 32725 29009 32759
rect 29009 32725 29043 32759
rect 29043 32725 29052 32759
rect 29000 32716 29052 32725
rect 29552 32759 29604 32768
rect 29552 32725 29561 32759
rect 29561 32725 29595 32759
rect 29595 32725 29604 32759
rect 29552 32716 29604 32725
rect 38752 32716 38804 32768
rect 41604 32716 41656 32768
rect 42616 32716 42668 32768
rect 44272 32716 44324 32768
rect 45192 32716 45244 32768
rect 47492 32852 47544 32904
rect 47860 32920 47912 32972
rect 50068 32920 50120 32972
rect 51816 32988 51868 33040
rect 57244 32988 57296 33040
rect 47952 32716 48004 32768
rect 49240 32784 49292 32836
rect 50160 32784 50212 32836
rect 49608 32716 49660 32768
rect 57152 32920 57204 32972
rect 57796 32963 57848 32972
rect 57796 32929 57805 32963
rect 57805 32929 57839 32963
rect 57839 32929 57848 32963
rect 57796 32920 57848 32929
rect 54116 32895 54168 32904
rect 50896 32827 50948 32836
rect 50896 32793 50905 32827
rect 50905 32793 50939 32827
rect 50939 32793 50948 32827
rect 50896 32784 50948 32793
rect 51080 32827 51132 32836
rect 51080 32793 51105 32827
rect 51105 32793 51132 32827
rect 51080 32784 51132 32793
rect 54116 32861 54125 32895
rect 54125 32861 54159 32895
rect 54159 32861 54168 32895
rect 54116 32852 54168 32861
rect 54576 32895 54628 32904
rect 54576 32861 54585 32895
rect 54585 32861 54619 32895
rect 54619 32861 54628 32895
rect 54576 32852 54628 32861
rect 54760 32895 54812 32904
rect 54760 32861 54769 32895
rect 54769 32861 54803 32895
rect 54803 32861 54812 32895
rect 54760 32852 54812 32861
rect 54208 32784 54260 32836
rect 55496 32827 55548 32836
rect 55496 32793 55505 32827
rect 55505 32793 55539 32827
rect 55539 32793 55548 32827
rect 55496 32784 55548 32793
rect 56600 32784 56652 32836
rect 53932 32716 53984 32768
rect 57152 32716 57204 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 25044 32512 25096 32564
rect 26240 32555 26292 32564
rect 26240 32521 26249 32555
rect 26249 32521 26283 32555
rect 26283 32521 26292 32555
rect 26240 32512 26292 32521
rect 40684 32512 40736 32564
rect 41604 32512 41656 32564
rect 42432 32555 42484 32564
rect 42432 32521 42441 32555
rect 42441 32521 42475 32555
rect 42475 32521 42484 32555
rect 42432 32512 42484 32521
rect 47400 32512 47452 32564
rect 24032 32419 24084 32428
rect 24032 32385 24041 32419
rect 24041 32385 24075 32419
rect 24075 32385 24084 32419
rect 24032 32376 24084 32385
rect 24952 32444 25004 32496
rect 25136 32419 25188 32428
rect 25136 32385 25170 32419
rect 25170 32385 25188 32419
rect 27160 32419 27212 32428
rect 25136 32376 25188 32385
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 29552 32376 29604 32428
rect 32312 32419 32364 32428
rect 32312 32385 32321 32419
rect 32321 32385 32355 32419
rect 32355 32385 32364 32419
rect 32312 32376 32364 32385
rect 34704 32444 34756 32496
rect 36728 32444 36780 32496
rect 41696 32444 41748 32496
rect 48320 32512 48372 32564
rect 48688 32487 48740 32496
rect 34796 32376 34848 32428
rect 35716 32376 35768 32428
rect 37188 32376 37240 32428
rect 41236 32419 41288 32428
rect 41236 32385 41245 32419
rect 41245 32385 41279 32419
rect 41279 32385 41288 32419
rect 41236 32376 41288 32385
rect 41512 32419 41564 32428
rect 41512 32385 41521 32419
rect 41521 32385 41555 32419
rect 41555 32385 41564 32419
rect 41512 32376 41564 32385
rect 41880 32376 41932 32428
rect 42248 32376 42300 32428
rect 42708 32419 42760 32428
rect 42708 32385 42717 32419
rect 42717 32385 42751 32419
rect 42751 32385 42760 32419
rect 42708 32376 42760 32385
rect 27620 32308 27672 32360
rect 30380 32308 30432 32360
rect 44456 32376 44508 32428
rect 45008 32419 45060 32428
rect 45008 32385 45017 32419
rect 45017 32385 45051 32419
rect 45051 32385 45060 32419
rect 45008 32376 45060 32385
rect 45192 32419 45244 32428
rect 45192 32385 45201 32419
rect 45201 32385 45235 32419
rect 45235 32385 45244 32419
rect 45192 32376 45244 32385
rect 43076 32308 43128 32360
rect 48044 32376 48096 32428
rect 48228 32419 48280 32428
rect 48228 32385 48237 32419
rect 48237 32385 48271 32419
rect 48271 32385 48280 32419
rect 48228 32376 48280 32385
rect 48688 32453 48697 32487
rect 48697 32453 48731 32487
rect 48731 32453 48740 32487
rect 48688 32444 48740 32453
rect 51540 32444 51592 32496
rect 51816 32487 51868 32496
rect 51816 32453 51825 32487
rect 51825 32453 51859 32487
rect 51859 32453 51868 32487
rect 51816 32444 51868 32453
rect 53748 32512 53800 32564
rect 56508 32555 56560 32564
rect 56508 32521 56517 32555
rect 56517 32521 56551 32555
rect 56551 32521 56560 32555
rect 56508 32512 56560 32521
rect 57060 32555 57112 32564
rect 57060 32521 57069 32555
rect 57069 32521 57103 32555
rect 57103 32521 57112 32555
rect 57060 32512 57112 32521
rect 48872 32419 48924 32428
rect 48872 32385 48881 32419
rect 48881 32385 48915 32419
rect 48915 32385 48924 32419
rect 48872 32376 48924 32385
rect 44456 32240 44508 32292
rect 47860 32240 47912 32292
rect 25228 32172 25280 32224
rect 25504 32172 25556 32224
rect 28724 32172 28776 32224
rect 31760 32172 31812 32224
rect 36728 32172 36780 32224
rect 38660 32215 38712 32224
rect 38660 32181 38669 32215
rect 38669 32181 38703 32215
rect 38703 32181 38712 32215
rect 38660 32172 38712 32181
rect 44824 32172 44876 32224
rect 50068 32376 50120 32428
rect 50896 32419 50948 32428
rect 50896 32385 50905 32419
rect 50905 32385 50939 32419
rect 50939 32385 50948 32419
rect 50896 32376 50948 32385
rect 51264 32376 51316 32428
rect 52644 32376 52696 32428
rect 53564 32376 53616 32428
rect 52552 32308 52604 32360
rect 53104 32308 53156 32360
rect 55496 32376 55548 32428
rect 56968 32419 57020 32428
rect 56968 32385 56977 32419
rect 56977 32385 57011 32419
rect 57011 32385 57020 32419
rect 56968 32376 57020 32385
rect 57152 32419 57204 32428
rect 57152 32385 57161 32419
rect 57161 32385 57195 32419
rect 57195 32385 57204 32419
rect 57152 32376 57204 32385
rect 55588 32308 55640 32360
rect 56600 32308 56652 32360
rect 49976 32240 50028 32292
rect 52828 32283 52880 32292
rect 52828 32249 52837 32283
rect 52837 32249 52871 32283
rect 52871 32249 52880 32283
rect 52828 32240 52880 32249
rect 54668 32240 54720 32292
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 28540 32011 28592 32020
rect 28540 31977 28549 32011
rect 28549 31977 28583 32011
rect 28583 31977 28592 32011
rect 28540 31968 28592 31977
rect 27988 31900 28040 31952
rect 25044 31875 25096 31884
rect 25044 31841 25053 31875
rect 25053 31841 25087 31875
rect 25087 31841 25096 31875
rect 25044 31832 25096 31841
rect 30380 31832 30432 31884
rect 26976 31764 27028 31816
rect 28724 31807 28776 31816
rect 28724 31773 28733 31807
rect 28733 31773 28767 31807
rect 28767 31773 28776 31807
rect 28724 31764 28776 31773
rect 30932 31832 30984 31884
rect 41420 31968 41472 32020
rect 42708 31968 42760 32020
rect 46940 31968 46992 32020
rect 38844 31900 38896 31952
rect 25504 31696 25556 31748
rect 33784 31832 33836 31884
rect 34704 31875 34756 31884
rect 34704 31841 34713 31875
rect 34713 31841 34747 31875
rect 34747 31841 34756 31875
rect 34704 31832 34756 31841
rect 37188 31875 37240 31884
rect 37188 31841 37197 31875
rect 37197 31841 37231 31875
rect 37231 31841 37240 31875
rect 37188 31832 37240 31841
rect 34520 31764 34572 31816
rect 37464 31807 37516 31816
rect 37464 31773 37498 31807
rect 37498 31773 37516 31807
rect 37464 31764 37516 31773
rect 43076 31900 43128 31952
rect 46756 31900 46808 31952
rect 42248 31807 42300 31816
rect 42248 31773 42257 31807
rect 42257 31773 42291 31807
rect 42291 31773 42300 31807
rect 42248 31764 42300 31773
rect 43444 31807 43496 31816
rect 43444 31773 43453 31807
rect 43453 31773 43487 31807
rect 43487 31773 43496 31807
rect 43444 31764 43496 31773
rect 43628 31807 43680 31816
rect 43628 31773 43637 31807
rect 43637 31773 43671 31807
rect 43671 31773 43680 31807
rect 43628 31764 43680 31773
rect 44272 31807 44324 31816
rect 44272 31773 44281 31807
rect 44281 31773 44315 31807
rect 44315 31773 44324 31807
rect 44272 31764 44324 31773
rect 44456 31807 44508 31816
rect 44456 31773 44465 31807
rect 44465 31773 44499 31807
rect 44499 31773 44508 31807
rect 44456 31764 44508 31773
rect 45192 31832 45244 31884
rect 46664 31832 46716 31884
rect 45008 31764 45060 31816
rect 46756 31764 46808 31816
rect 34704 31696 34756 31748
rect 35808 31696 35860 31748
rect 48688 31968 48740 32020
rect 48872 32011 48924 32020
rect 48872 31977 48881 32011
rect 48881 31977 48915 32011
rect 48915 31977 48924 32011
rect 48872 31968 48924 31977
rect 53104 31968 53156 32020
rect 53564 32011 53616 32020
rect 53564 31977 53573 32011
rect 53573 31977 53607 32011
rect 53607 31977 53616 32011
rect 53564 31968 53616 31977
rect 55404 31968 55456 32020
rect 48320 31900 48372 31952
rect 49424 31900 49476 31952
rect 54760 31900 54812 31952
rect 56048 31900 56100 31952
rect 52828 31832 52880 31884
rect 47952 31807 48004 31816
rect 47952 31773 47961 31807
rect 47961 31773 47995 31807
rect 47995 31773 48004 31807
rect 47952 31764 48004 31773
rect 50896 31807 50948 31816
rect 50896 31773 50905 31807
rect 50905 31773 50939 31807
rect 50939 31773 50948 31807
rect 50896 31764 50948 31773
rect 51080 31764 51132 31816
rect 49976 31696 50028 31748
rect 32496 31671 32548 31680
rect 32496 31637 32505 31671
rect 32505 31637 32539 31671
rect 32539 31637 32548 31671
rect 32496 31628 32548 31637
rect 34980 31628 35032 31680
rect 35716 31628 35768 31680
rect 47124 31628 47176 31680
rect 47308 31628 47360 31680
rect 51356 31628 51408 31680
rect 52552 31764 52604 31816
rect 52644 31807 52696 31816
rect 52644 31773 52653 31807
rect 52653 31773 52687 31807
rect 52687 31773 52696 31807
rect 52644 31764 52696 31773
rect 53472 31764 53524 31816
rect 53748 31764 53800 31816
rect 55864 31807 55916 31816
rect 55864 31773 55873 31807
rect 55873 31773 55907 31807
rect 55907 31773 55916 31807
rect 55864 31764 55916 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 25136 31424 25188 31476
rect 29000 31424 29052 31476
rect 30932 31424 30984 31476
rect 26240 31356 26292 31408
rect 25228 31331 25280 31340
rect 25228 31297 25237 31331
rect 25237 31297 25271 31331
rect 25271 31297 25280 31331
rect 25228 31288 25280 31297
rect 27620 31288 27672 31340
rect 28172 31288 28224 31340
rect 31760 31356 31812 31408
rect 31852 31356 31904 31408
rect 31116 31288 31168 31340
rect 32220 31288 32272 31340
rect 32496 31331 32548 31340
rect 32496 31297 32505 31331
rect 32505 31297 32539 31331
rect 32539 31297 32548 31331
rect 32496 31288 32548 31297
rect 34704 31288 34756 31340
rect 34980 31331 35032 31340
rect 34980 31297 34989 31331
rect 34989 31297 35023 31331
rect 35023 31297 35032 31331
rect 34980 31288 35032 31297
rect 35900 31424 35952 31476
rect 39212 31424 39264 31476
rect 39672 31424 39724 31476
rect 40316 31424 40368 31476
rect 43076 31424 43128 31476
rect 43628 31424 43680 31476
rect 37648 31356 37700 31408
rect 35808 31288 35860 31340
rect 38660 31288 38712 31340
rect 39396 31288 39448 31340
rect 41512 31356 41564 31408
rect 28816 31220 28868 31272
rect 30288 31220 30340 31272
rect 39120 31152 39172 31204
rect 40960 31288 41012 31340
rect 43536 31288 43588 31340
rect 45284 31424 45336 31476
rect 46480 31424 46532 31476
rect 48136 31467 48188 31476
rect 48136 31433 48145 31467
rect 48145 31433 48179 31467
rect 48179 31433 48188 31467
rect 48136 31424 48188 31433
rect 49700 31467 49752 31476
rect 49700 31433 49709 31467
rect 49709 31433 49743 31467
rect 49743 31433 49752 31467
rect 49700 31424 49752 31433
rect 51264 31424 51316 31476
rect 49240 31356 49292 31408
rect 44824 31331 44876 31340
rect 44824 31297 44833 31331
rect 44833 31297 44867 31331
rect 44867 31297 44876 31331
rect 44824 31288 44876 31297
rect 46112 31331 46164 31340
rect 46112 31297 46121 31331
rect 46121 31297 46155 31331
rect 46155 31297 46164 31331
rect 46112 31288 46164 31297
rect 47584 31331 47636 31340
rect 47584 31297 47593 31331
rect 47593 31297 47627 31331
rect 47627 31297 47636 31331
rect 47584 31288 47636 31297
rect 44272 31220 44324 31272
rect 44456 31220 44508 31272
rect 43444 31152 43496 31204
rect 45284 31220 45336 31272
rect 48044 31288 48096 31340
rect 49332 31331 49384 31340
rect 49332 31297 49341 31331
rect 49341 31297 49375 31331
rect 49375 31297 49384 31331
rect 49332 31288 49384 31297
rect 49240 31220 49292 31272
rect 49516 31331 49568 31340
rect 49516 31297 49525 31331
rect 49525 31297 49559 31331
rect 49559 31297 49568 31331
rect 50712 31356 50764 31408
rect 51172 31399 51224 31408
rect 51172 31365 51181 31399
rect 51181 31365 51215 31399
rect 51215 31365 51224 31399
rect 51172 31356 51224 31365
rect 53012 31424 53064 31476
rect 54576 31424 54628 31476
rect 52184 31356 52236 31408
rect 53748 31399 53800 31408
rect 53748 31365 53757 31399
rect 53757 31365 53791 31399
rect 53791 31365 53800 31399
rect 53748 31356 53800 31365
rect 49516 31288 49568 31297
rect 50896 31288 50948 31340
rect 51080 31331 51132 31340
rect 51080 31297 51089 31331
rect 51089 31297 51123 31331
rect 51123 31297 51132 31331
rect 52000 31331 52052 31340
rect 51080 31288 51132 31297
rect 49976 31220 50028 31272
rect 52000 31297 52009 31331
rect 52009 31297 52043 31331
rect 52043 31297 52052 31331
rect 52000 31288 52052 31297
rect 52368 31288 52420 31340
rect 53472 31331 53524 31340
rect 27712 31084 27764 31136
rect 29000 31084 29052 31136
rect 30196 31127 30248 31136
rect 30196 31093 30205 31127
rect 30205 31093 30239 31127
rect 30239 31093 30248 31127
rect 30196 31084 30248 31093
rect 32312 31084 32364 31136
rect 36636 31084 36688 31136
rect 38844 31084 38896 31136
rect 39028 31084 39080 31136
rect 39488 31127 39540 31136
rect 39488 31093 39497 31127
rect 39497 31093 39531 31127
rect 39531 31093 39540 31127
rect 39488 31084 39540 31093
rect 44180 31127 44232 31136
rect 44180 31093 44189 31127
rect 44189 31093 44223 31127
rect 44223 31093 44232 31127
rect 44180 31084 44232 31093
rect 44364 31084 44416 31136
rect 44732 31084 44784 31136
rect 51908 31152 51960 31204
rect 52828 31152 52880 31204
rect 48228 31084 48280 31136
rect 51172 31084 51224 31136
rect 53472 31297 53481 31331
rect 53481 31297 53515 31331
rect 53515 31297 53524 31331
rect 53472 31288 53524 31297
rect 53564 31331 53616 31340
rect 53564 31297 53573 31331
rect 53573 31297 53607 31331
rect 53607 31297 53616 31331
rect 55404 31424 55456 31476
rect 55588 31467 55640 31476
rect 55588 31433 55597 31467
rect 55597 31433 55631 31467
rect 55631 31433 55640 31467
rect 55588 31424 55640 31433
rect 56140 31424 56192 31476
rect 56600 31467 56652 31476
rect 56600 31433 56609 31467
rect 56609 31433 56643 31467
rect 56643 31433 56652 31467
rect 56600 31424 56652 31433
rect 55864 31356 55916 31408
rect 53564 31288 53616 31297
rect 55772 31331 55824 31340
rect 53656 31152 53708 31204
rect 55772 31297 55781 31331
rect 55781 31297 55815 31331
rect 55815 31297 55824 31331
rect 55772 31288 55824 31297
rect 56048 31331 56100 31340
rect 56048 31297 56057 31331
rect 56057 31297 56091 31331
rect 56091 31297 56100 31331
rect 56048 31288 56100 31297
rect 55588 31152 55640 31204
rect 56140 31152 56192 31204
rect 56324 31084 56376 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 28172 30880 28224 30932
rect 31208 30880 31260 30932
rect 36728 30923 36780 30932
rect 36728 30889 36737 30923
rect 36737 30889 36771 30923
rect 36771 30889 36780 30923
rect 36728 30880 36780 30889
rect 39028 30923 39080 30932
rect 39028 30889 39037 30923
rect 39037 30889 39071 30923
rect 39071 30889 39080 30923
rect 39028 30880 39080 30889
rect 44824 30880 44876 30932
rect 46296 30923 46348 30932
rect 46296 30889 46305 30923
rect 46305 30889 46339 30923
rect 46339 30889 46348 30923
rect 46296 30880 46348 30889
rect 47952 30880 48004 30932
rect 49148 30923 49200 30932
rect 49148 30889 49157 30923
rect 49157 30889 49191 30923
rect 49191 30889 49200 30923
rect 49148 30880 49200 30889
rect 50712 30923 50764 30932
rect 50712 30889 50721 30923
rect 50721 30889 50755 30923
rect 50755 30889 50764 30923
rect 50712 30880 50764 30889
rect 51356 30923 51408 30932
rect 51356 30889 51365 30923
rect 51365 30889 51399 30923
rect 51399 30889 51408 30923
rect 51356 30880 51408 30889
rect 39396 30812 39448 30864
rect 41328 30812 41380 30864
rect 48780 30812 48832 30864
rect 30288 30744 30340 30796
rect 38936 30787 38988 30796
rect 38936 30753 38945 30787
rect 38945 30753 38979 30787
rect 38979 30753 38988 30787
rect 38936 30744 38988 30753
rect 27712 30719 27764 30728
rect 27712 30685 27721 30719
rect 27721 30685 27755 30719
rect 27755 30685 27764 30719
rect 27712 30676 27764 30685
rect 29276 30676 29328 30728
rect 34704 30676 34756 30728
rect 35532 30676 35584 30728
rect 36636 30719 36688 30728
rect 36636 30685 36645 30719
rect 36645 30685 36679 30719
rect 36679 30685 36688 30719
rect 36636 30676 36688 30685
rect 36728 30676 36780 30728
rect 41512 30744 41564 30796
rect 39120 30719 39172 30728
rect 39120 30685 39129 30719
rect 39129 30685 39163 30719
rect 39163 30685 39172 30719
rect 39120 30676 39172 30685
rect 39304 30676 39356 30728
rect 39948 30719 40000 30728
rect 39948 30685 39957 30719
rect 39957 30685 39991 30719
rect 39991 30685 40000 30719
rect 39948 30676 40000 30685
rect 43444 30719 43496 30728
rect 30196 30608 30248 30660
rect 37188 30608 37240 30660
rect 27528 30583 27580 30592
rect 27528 30549 27537 30583
rect 27537 30549 27571 30583
rect 27571 30549 27580 30583
rect 27528 30540 27580 30549
rect 28356 30540 28408 30592
rect 37096 30583 37148 30592
rect 37096 30549 37105 30583
rect 37105 30549 37139 30583
rect 37139 30549 37148 30583
rect 37096 30540 37148 30549
rect 40408 30608 40460 30660
rect 43444 30685 43453 30719
rect 43453 30685 43487 30719
rect 43487 30685 43496 30719
rect 43444 30676 43496 30685
rect 44548 30744 44600 30796
rect 45284 30787 45336 30796
rect 45284 30753 45293 30787
rect 45293 30753 45327 30787
rect 45327 30753 45336 30787
rect 45284 30744 45336 30753
rect 44272 30719 44324 30728
rect 44272 30685 44281 30719
rect 44281 30685 44315 30719
rect 44315 30685 44324 30719
rect 44272 30676 44324 30685
rect 46480 30719 46532 30728
rect 46480 30685 46489 30719
rect 46489 30685 46523 30719
rect 46523 30685 46532 30719
rect 46480 30676 46532 30685
rect 46756 30719 46808 30728
rect 46756 30685 46765 30719
rect 46765 30685 46799 30719
rect 46799 30685 46808 30719
rect 46756 30676 46808 30685
rect 47124 30676 47176 30728
rect 51080 30744 51132 30796
rect 48872 30719 48924 30728
rect 48872 30685 48881 30719
rect 48881 30685 48915 30719
rect 48915 30685 48924 30719
rect 48872 30676 48924 30685
rect 49700 30676 49752 30728
rect 51172 30676 51224 30728
rect 52644 30880 52696 30932
rect 56048 30880 56100 30932
rect 56324 30787 56376 30796
rect 56324 30753 56333 30787
rect 56333 30753 56367 30787
rect 56367 30753 56376 30787
rect 56324 30744 56376 30753
rect 44364 30608 44416 30660
rect 40224 30540 40276 30592
rect 40592 30540 40644 30592
rect 41328 30583 41380 30592
rect 41328 30549 41337 30583
rect 41337 30549 41371 30583
rect 41371 30549 41380 30583
rect 41328 30540 41380 30549
rect 43536 30583 43588 30592
rect 43536 30549 43545 30583
rect 43545 30549 43579 30583
rect 43579 30549 43588 30583
rect 43536 30540 43588 30549
rect 44732 30608 44784 30660
rect 47768 30608 47820 30660
rect 50988 30608 51040 30660
rect 54668 30719 54720 30728
rect 52092 30651 52144 30660
rect 52092 30617 52101 30651
rect 52101 30617 52135 30651
rect 52135 30617 52144 30651
rect 52092 30608 52144 30617
rect 52368 30608 52420 30660
rect 54668 30685 54677 30719
rect 54677 30685 54711 30719
rect 54711 30685 54720 30719
rect 54668 30676 54720 30685
rect 55588 30719 55640 30728
rect 55588 30685 55597 30719
rect 55597 30685 55631 30719
rect 55631 30685 55640 30719
rect 55588 30676 55640 30685
rect 54760 30608 54812 30660
rect 55404 30651 55456 30660
rect 55404 30617 55413 30651
rect 55413 30617 55447 30651
rect 55447 30617 55456 30651
rect 55404 30608 55456 30617
rect 57980 30608 58032 30660
rect 58164 30651 58216 30660
rect 58164 30617 58173 30651
rect 58173 30617 58207 30651
rect 58207 30617 58216 30651
rect 58164 30608 58216 30617
rect 46572 30540 46624 30592
rect 50160 30540 50212 30592
rect 54208 30540 54260 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 28356 30379 28408 30388
rect 28356 30345 28365 30379
rect 28365 30345 28399 30379
rect 28399 30345 28408 30379
rect 28356 30336 28408 30345
rect 35532 30336 35584 30388
rect 38660 30379 38712 30388
rect 27528 30268 27580 30320
rect 34152 30311 34204 30320
rect 34152 30277 34186 30311
rect 34186 30277 34204 30311
rect 38660 30345 38669 30379
rect 38669 30345 38703 30379
rect 38703 30345 38712 30379
rect 38660 30336 38712 30345
rect 38844 30336 38896 30388
rect 40316 30379 40368 30388
rect 34152 30268 34204 30277
rect 2412 30243 2464 30252
rect 2412 30209 2421 30243
rect 2421 30209 2455 30243
rect 2455 30209 2464 30243
rect 2412 30200 2464 30209
rect 24584 30200 24636 30252
rect 26976 30243 27028 30252
rect 26976 30209 26985 30243
rect 26985 30209 27019 30243
rect 27019 30209 27028 30243
rect 26976 30200 27028 30209
rect 28080 30200 28132 30252
rect 28816 30200 28868 30252
rect 31116 30175 31168 30184
rect 1952 30039 2004 30048
rect 1952 30005 1961 30039
rect 1961 30005 1995 30039
rect 1995 30005 2004 30039
rect 1952 29996 2004 30005
rect 2136 29996 2188 30048
rect 26056 30039 26108 30048
rect 26056 30005 26065 30039
rect 26065 30005 26099 30039
rect 26099 30005 26108 30039
rect 26056 29996 26108 30005
rect 31116 30141 31125 30175
rect 31125 30141 31159 30175
rect 31159 30141 31168 30175
rect 31116 30132 31168 30141
rect 33784 30200 33836 30252
rect 37096 30268 37148 30320
rect 31944 30132 31996 30184
rect 38660 30200 38712 30252
rect 40316 30345 40325 30379
rect 40325 30345 40359 30379
rect 40359 30345 40368 30379
rect 40316 30336 40368 30345
rect 43444 30336 43496 30388
rect 41880 30311 41932 30320
rect 41880 30277 41889 30311
rect 41889 30277 41923 30311
rect 41923 30277 41932 30311
rect 41880 30268 41932 30277
rect 43536 30268 43588 30320
rect 39948 30243 40000 30252
rect 39948 30209 39957 30243
rect 39957 30209 39991 30243
rect 39991 30209 40000 30243
rect 39948 30200 40000 30209
rect 31668 30064 31720 30116
rect 38568 30132 38620 30184
rect 40500 30132 40552 30184
rect 29092 30039 29144 30048
rect 29092 30005 29101 30039
rect 29101 30005 29135 30039
rect 29135 30005 29144 30039
rect 29092 29996 29144 30005
rect 30472 29996 30524 30048
rect 30840 29996 30892 30048
rect 35808 29996 35860 30048
rect 36452 30039 36504 30048
rect 36452 30005 36461 30039
rect 36461 30005 36495 30039
rect 36495 30005 36504 30039
rect 36452 29996 36504 30005
rect 37648 30039 37700 30048
rect 37648 30005 37657 30039
rect 37657 30005 37691 30039
rect 37691 30005 37700 30039
rect 37648 29996 37700 30005
rect 37740 29996 37792 30048
rect 40316 30039 40368 30048
rect 40316 30005 40325 30039
rect 40325 30005 40359 30039
rect 40359 30005 40368 30039
rect 40316 29996 40368 30005
rect 40500 30039 40552 30048
rect 40500 30005 40509 30039
rect 40509 30005 40543 30039
rect 40543 30005 40552 30039
rect 40500 29996 40552 30005
rect 41604 30200 41656 30252
rect 42432 30243 42484 30252
rect 42432 30209 42441 30243
rect 42441 30209 42475 30243
rect 42475 30209 42484 30243
rect 42432 30200 42484 30209
rect 42708 30200 42760 30252
rect 43996 30200 44048 30252
rect 44548 30336 44600 30388
rect 45468 30336 45520 30388
rect 49148 30336 49200 30388
rect 55772 30379 55824 30388
rect 55772 30345 55781 30379
rect 55781 30345 55815 30379
rect 55815 30345 55824 30379
rect 55772 30336 55824 30345
rect 44916 30268 44968 30320
rect 49332 30268 49384 30320
rect 42064 30132 42116 30184
rect 43352 30132 43404 30184
rect 43812 30132 43864 30184
rect 43536 30064 43588 30116
rect 45192 30243 45244 30252
rect 44916 30132 44968 30184
rect 45192 30209 45201 30243
rect 45201 30209 45235 30243
rect 45235 30209 45244 30243
rect 45192 30200 45244 30209
rect 46756 30200 46808 30252
rect 47952 30200 48004 30252
rect 45100 30132 45152 30184
rect 48688 30200 48740 30252
rect 49240 30200 49292 30252
rect 50988 30268 51040 30320
rect 54208 30268 54260 30320
rect 57980 30311 58032 30320
rect 57980 30277 57989 30311
rect 57989 30277 58023 30311
rect 58023 30277 58032 30311
rect 57980 30268 58032 30277
rect 49516 30200 49568 30252
rect 51264 30200 51316 30252
rect 52092 30200 52144 30252
rect 54668 30243 54720 30252
rect 54668 30209 54677 30243
rect 54677 30209 54711 30243
rect 54711 30209 54720 30243
rect 54668 30200 54720 30209
rect 54760 30243 54812 30252
rect 54760 30209 54769 30243
rect 54769 30209 54803 30243
rect 54803 30209 54812 30243
rect 54760 30200 54812 30209
rect 56692 30200 56744 30252
rect 57336 30200 57388 30252
rect 57612 30200 57664 30252
rect 49976 30132 50028 30184
rect 50804 30175 50856 30184
rect 50804 30141 50813 30175
rect 50813 30141 50847 30175
rect 50847 30141 50856 30175
rect 50804 30132 50856 30141
rect 49516 30064 49568 30116
rect 49608 30064 49660 30116
rect 52000 30064 52052 30116
rect 48136 30039 48188 30048
rect 48136 30005 48145 30039
rect 48145 30005 48179 30039
rect 48179 30005 48188 30039
rect 48136 29996 48188 30005
rect 56508 29996 56560 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 31852 29792 31904 29844
rect 38660 29792 38712 29844
rect 38752 29792 38804 29844
rect 39764 29792 39816 29844
rect 42248 29792 42300 29844
rect 45192 29792 45244 29844
rect 24584 29588 24636 29640
rect 30840 29724 30892 29776
rect 36452 29724 36504 29776
rect 40040 29724 40092 29776
rect 40224 29767 40276 29776
rect 40224 29733 40233 29767
rect 40233 29733 40267 29767
rect 40267 29733 40276 29767
rect 40224 29724 40276 29733
rect 40408 29724 40460 29776
rect 43536 29724 43588 29776
rect 27988 29699 28040 29708
rect 27988 29665 27997 29699
rect 27997 29665 28031 29699
rect 28031 29665 28040 29699
rect 27988 29656 28040 29665
rect 28080 29699 28132 29708
rect 28080 29665 28089 29699
rect 28089 29665 28123 29699
rect 28123 29665 28132 29699
rect 28080 29656 28132 29665
rect 31116 29656 31168 29708
rect 31944 29699 31996 29708
rect 28356 29588 28408 29640
rect 30840 29631 30892 29640
rect 27344 29520 27396 29572
rect 30840 29597 30849 29631
rect 30849 29597 30883 29631
rect 30883 29597 30892 29631
rect 30840 29588 30892 29597
rect 31944 29665 31953 29699
rect 31953 29665 31987 29699
rect 31987 29665 31996 29699
rect 31944 29656 31996 29665
rect 30472 29520 30524 29572
rect 33140 29588 33192 29640
rect 36636 29656 36688 29708
rect 38476 29656 38528 29708
rect 40500 29656 40552 29708
rect 42616 29656 42668 29708
rect 43444 29656 43496 29708
rect 37004 29631 37056 29640
rect 37004 29597 37013 29631
rect 37013 29597 37047 29631
rect 37047 29597 37056 29631
rect 37004 29588 37056 29597
rect 37188 29588 37240 29640
rect 38752 29631 38804 29640
rect 38752 29597 38761 29631
rect 38761 29597 38795 29631
rect 38795 29597 38804 29631
rect 38752 29588 38804 29597
rect 31760 29520 31812 29572
rect 32496 29520 32548 29572
rect 33692 29563 33744 29572
rect 33692 29529 33701 29563
rect 33701 29529 33735 29563
rect 33735 29529 33744 29563
rect 33692 29520 33744 29529
rect 28540 29452 28592 29504
rect 31944 29495 31996 29504
rect 31944 29461 31953 29495
rect 31953 29461 31987 29495
rect 31987 29461 31996 29495
rect 31944 29452 31996 29461
rect 36268 29452 36320 29504
rect 39580 29520 39632 29572
rect 40132 29631 40184 29640
rect 40132 29597 40141 29631
rect 40141 29597 40175 29631
rect 40175 29597 40184 29631
rect 40132 29588 40184 29597
rect 40408 29588 40460 29640
rect 40960 29631 41012 29640
rect 40960 29597 40969 29631
rect 40969 29597 41003 29631
rect 41003 29597 41012 29631
rect 40960 29588 41012 29597
rect 42064 29631 42116 29640
rect 42064 29597 42073 29631
rect 42073 29597 42107 29631
rect 42107 29597 42116 29631
rect 42064 29588 42116 29597
rect 43812 29631 43864 29640
rect 40224 29520 40276 29572
rect 43168 29520 43220 29572
rect 43812 29597 43821 29631
rect 43821 29597 43855 29631
rect 43855 29597 43864 29631
rect 43812 29588 43864 29597
rect 43996 29631 44048 29640
rect 43996 29597 44005 29631
rect 44005 29597 44039 29631
rect 44039 29597 44048 29631
rect 43996 29588 44048 29597
rect 44180 29588 44232 29640
rect 44916 29588 44968 29640
rect 43720 29563 43772 29572
rect 43720 29529 43729 29563
rect 43729 29529 43763 29563
rect 43763 29529 43772 29563
rect 46388 29792 46440 29844
rect 47584 29792 47636 29844
rect 52736 29792 52788 29844
rect 54024 29835 54076 29844
rect 54024 29801 54033 29835
rect 54033 29801 54067 29835
rect 54067 29801 54076 29835
rect 54024 29792 54076 29801
rect 55404 29835 55456 29844
rect 55404 29801 55413 29835
rect 55413 29801 55447 29835
rect 55447 29801 55456 29835
rect 55404 29792 55456 29801
rect 46756 29724 46808 29776
rect 47860 29724 47912 29776
rect 50160 29724 50212 29776
rect 48780 29656 48832 29708
rect 47584 29631 47636 29640
rect 47584 29597 47593 29631
rect 47593 29597 47627 29631
rect 47627 29597 47636 29631
rect 47584 29588 47636 29597
rect 48136 29588 48188 29640
rect 51172 29588 51224 29640
rect 51448 29631 51500 29640
rect 51448 29597 51457 29631
rect 51457 29597 51491 29631
rect 51491 29597 51500 29631
rect 51448 29588 51500 29597
rect 54024 29656 54076 29708
rect 56508 29699 56560 29708
rect 54208 29631 54260 29640
rect 46572 29563 46624 29572
rect 43720 29520 43772 29529
rect 46572 29529 46581 29563
rect 46581 29529 46615 29563
rect 46615 29529 46624 29563
rect 46572 29520 46624 29529
rect 47768 29520 47820 29572
rect 54208 29597 54217 29631
rect 54217 29597 54251 29631
rect 54251 29597 54260 29631
rect 54208 29588 54260 29597
rect 56508 29665 56517 29699
rect 56517 29665 56551 29699
rect 56551 29665 56560 29699
rect 56508 29656 56560 29665
rect 57888 29699 57940 29708
rect 57888 29665 57897 29699
rect 57897 29665 57931 29699
rect 57931 29665 57940 29699
rect 57888 29656 57940 29665
rect 55312 29631 55364 29640
rect 55312 29597 55321 29631
rect 55321 29597 55355 29631
rect 55355 29597 55364 29631
rect 55312 29588 55364 29597
rect 55496 29631 55548 29640
rect 55496 29597 55505 29631
rect 55505 29597 55539 29631
rect 55539 29597 55548 29631
rect 55496 29588 55548 29597
rect 56140 29588 56192 29640
rect 56324 29631 56376 29640
rect 56324 29597 56333 29631
rect 56333 29597 56367 29631
rect 56367 29597 56376 29631
rect 56324 29588 56376 29597
rect 52460 29520 52512 29572
rect 39212 29452 39264 29504
rect 39304 29452 39356 29504
rect 41052 29495 41104 29504
rect 41052 29461 41061 29495
rect 41061 29461 41095 29495
rect 41095 29461 41104 29495
rect 41052 29452 41104 29461
rect 43536 29452 43588 29504
rect 49884 29452 49936 29504
rect 53012 29452 53064 29504
rect 54392 29495 54444 29504
rect 54392 29461 54401 29495
rect 54401 29461 54435 29495
rect 54435 29461 54444 29495
rect 54392 29452 54444 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 28080 29248 28132 29300
rect 42616 29291 42668 29300
rect 2136 29223 2188 29232
rect 2136 29189 2145 29223
rect 2145 29189 2179 29223
rect 2179 29189 2188 29223
rect 2136 29180 2188 29189
rect 1952 29155 2004 29164
rect 1952 29121 1961 29155
rect 1961 29121 1995 29155
rect 1995 29121 2004 29155
rect 1952 29112 2004 29121
rect 24584 29155 24636 29164
rect 24584 29121 24593 29155
rect 24593 29121 24627 29155
rect 24627 29121 24636 29155
rect 24584 29112 24636 29121
rect 26976 29155 27028 29164
rect 26976 29121 26985 29155
rect 26985 29121 27019 29155
rect 27019 29121 27028 29155
rect 26976 29112 27028 29121
rect 27252 29155 27304 29164
rect 27252 29121 27286 29155
rect 27286 29121 27304 29155
rect 27252 29112 27304 29121
rect 30472 29112 30524 29164
rect 31024 29112 31076 29164
rect 37924 29112 37976 29164
rect 38476 29155 38528 29164
rect 38476 29121 38485 29155
rect 38485 29121 38519 29155
rect 38519 29121 38528 29155
rect 38476 29112 38528 29121
rect 2780 29087 2832 29096
rect 2780 29053 2789 29087
rect 2789 29053 2823 29087
rect 2823 29053 2832 29087
rect 2780 29044 2832 29053
rect 25228 29044 25280 29096
rect 3424 28976 3476 29028
rect 31760 29044 31812 29096
rect 32220 29087 32272 29096
rect 32220 29053 32229 29087
rect 32229 29053 32263 29087
rect 32263 29053 32272 29087
rect 32220 29044 32272 29053
rect 37372 29087 37424 29096
rect 37372 29053 37381 29087
rect 37381 29053 37415 29087
rect 37415 29053 37424 29087
rect 37372 29044 37424 29053
rect 30840 28976 30892 29028
rect 33508 29019 33560 29028
rect 33508 28985 33517 29019
rect 33517 28985 33551 29019
rect 33551 28985 33560 29019
rect 33508 28976 33560 28985
rect 36728 28976 36780 29028
rect 37004 28976 37056 29028
rect 38844 29155 38896 29164
rect 38844 29121 38853 29155
rect 38853 29121 38887 29155
rect 38887 29121 38896 29155
rect 38844 29112 38896 29121
rect 42616 29257 42625 29291
rect 42625 29257 42659 29291
rect 42659 29257 42668 29291
rect 42616 29248 42668 29257
rect 43352 29291 43404 29300
rect 43352 29257 43361 29291
rect 43361 29257 43395 29291
rect 43395 29257 43404 29291
rect 43352 29248 43404 29257
rect 44272 29248 44324 29300
rect 49976 29291 50028 29300
rect 49976 29257 49985 29291
rect 49985 29257 50019 29291
rect 50019 29257 50028 29291
rect 49976 29248 50028 29257
rect 50620 29248 50672 29300
rect 50988 29291 51040 29300
rect 50988 29257 50997 29291
rect 50997 29257 51031 29291
rect 51031 29257 51040 29291
rect 51816 29291 51868 29300
rect 50988 29248 51040 29257
rect 51816 29257 51825 29291
rect 51825 29257 51859 29291
rect 51859 29257 51868 29291
rect 51816 29248 51868 29257
rect 39580 29180 39632 29232
rect 43444 29180 43496 29232
rect 48688 29180 48740 29232
rect 49424 29180 49476 29232
rect 40592 29112 40644 29164
rect 40960 29112 41012 29164
rect 42432 29112 42484 29164
rect 42708 29155 42760 29164
rect 42708 29121 42717 29155
rect 42717 29121 42751 29155
rect 42751 29121 42760 29155
rect 42708 29112 42760 29121
rect 43168 29155 43220 29164
rect 43168 29121 43177 29155
rect 43177 29121 43211 29155
rect 43211 29121 43220 29155
rect 43168 29112 43220 29121
rect 44180 29112 44232 29164
rect 38660 28976 38712 29028
rect 41144 28976 41196 29028
rect 43996 29044 44048 29096
rect 46664 29112 46716 29164
rect 49792 29112 49844 29164
rect 49884 29155 49936 29164
rect 49884 29121 49893 29155
rect 49893 29121 49927 29155
rect 49927 29121 49936 29155
rect 49884 29112 49936 29121
rect 52460 29180 52512 29232
rect 46480 29044 46532 29096
rect 50068 29044 50120 29096
rect 50988 29044 51040 29096
rect 45652 28976 45704 29028
rect 50620 28976 50672 29028
rect 51448 29112 51500 29164
rect 54392 29248 54444 29300
rect 54760 29248 54812 29300
rect 52920 29087 52972 29096
rect 52920 29053 52929 29087
rect 52929 29053 52963 29087
rect 52963 29053 52972 29087
rect 52920 29044 52972 29053
rect 53012 29087 53064 29096
rect 53012 29053 53021 29087
rect 53021 29053 53055 29087
rect 53055 29053 53064 29087
rect 53012 29044 53064 29053
rect 54024 29087 54076 29096
rect 52828 28976 52880 29028
rect 54024 29053 54033 29087
rect 54033 29053 54067 29087
rect 54067 29053 54076 29087
rect 54024 29044 54076 29053
rect 31484 28908 31536 28960
rect 32312 28951 32364 28960
rect 32312 28917 32321 28951
rect 32321 28917 32355 28951
rect 32355 28917 32364 28951
rect 32312 28908 32364 28917
rect 37464 28951 37516 28960
rect 37464 28917 37473 28951
rect 37473 28917 37507 28951
rect 37507 28917 37516 28951
rect 37464 28908 37516 28917
rect 38016 28908 38068 28960
rect 38292 28951 38344 28960
rect 38292 28917 38301 28951
rect 38301 28917 38335 28951
rect 38335 28917 38344 28951
rect 38292 28908 38344 28917
rect 40868 28908 40920 28960
rect 42524 28908 42576 28960
rect 45928 28951 45980 28960
rect 45928 28917 45937 28951
rect 45937 28917 45971 28951
rect 45971 28917 45980 28951
rect 45928 28908 45980 28917
rect 46020 28908 46072 28960
rect 48504 28908 48556 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 25228 28747 25280 28756
rect 25228 28713 25237 28747
rect 25237 28713 25271 28747
rect 25271 28713 25280 28747
rect 25228 28704 25280 28713
rect 27252 28704 27304 28756
rect 28264 28704 28316 28756
rect 40868 28704 40920 28756
rect 28540 28611 28592 28620
rect 28540 28577 28549 28611
rect 28549 28577 28583 28611
rect 28583 28577 28592 28611
rect 28540 28568 28592 28577
rect 24860 28364 24912 28416
rect 26148 28500 26200 28552
rect 27160 28543 27212 28552
rect 27160 28509 27169 28543
rect 27169 28509 27203 28543
rect 27203 28509 27212 28543
rect 27160 28500 27212 28509
rect 27344 28543 27396 28552
rect 27344 28509 27353 28543
rect 27353 28509 27387 28543
rect 27387 28509 27396 28543
rect 27344 28500 27396 28509
rect 32312 28636 32364 28688
rect 29000 28500 29052 28552
rect 31944 28568 31996 28620
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 29828 28500 29880 28509
rect 31116 28500 31168 28552
rect 32680 28543 32732 28552
rect 32680 28509 32689 28543
rect 32689 28509 32723 28543
rect 32723 28509 32732 28543
rect 32680 28500 32732 28509
rect 32864 28543 32916 28552
rect 32864 28509 32873 28543
rect 32873 28509 32907 28543
rect 32907 28509 32916 28543
rect 32864 28500 32916 28509
rect 30380 28432 30432 28484
rect 36820 28636 36872 28688
rect 34704 28611 34756 28620
rect 34704 28577 34713 28611
rect 34713 28577 34747 28611
rect 34747 28577 34756 28611
rect 34704 28568 34756 28577
rect 35808 28568 35860 28620
rect 40776 28636 40828 28688
rect 47492 28704 47544 28756
rect 47952 28704 48004 28756
rect 48780 28747 48832 28756
rect 48780 28713 48789 28747
rect 48789 28713 48823 28747
rect 48823 28713 48832 28747
rect 48780 28704 48832 28713
rect 52828 28747 52880 28756
rect 52828 28713 52837 28747
rect 52837 28713 52871 28747
rect 52871 28713 52880 28747
rect 52828 28704 52880 28713
rect 53012 28704 53064 28756
rect 55312 28704 55364 28756
rect 42524 28636 42576 28688
rect 55220 28636 55272 28688
rect 37740 28543 37792 28552
rect 37740 28509 37749 28543
rect 37749 28509 37783 28543
rect 37783 28509 37792 28543
rect 37740 28500 37792 28509
rect 38016 28543 38068 28552
rect 38016 28509 38025 28543
rect 38025 28509 38059 28543
rect 38059 28509 38068 28543
rect 38016 28500 38068 28509
rect 38936 28500 38988 28552
rect 35624 28432 35676 28484
rect 37188 28432 37240 28484
rect 37280 28432 37332 28484
rect 40960 28500 41012 28552
rect 41144 28543 41196 28552
rect 41144 28509 41153 28543
rect 41153 28509 41187 28543
rect 41187 28509 41196 28543
rect 41144 28500 41196 28509
rect 42892 28568 42944 28620
rect 43352 28568 43404 28620
rect 41788 28500 41840 28552
rect 43720 28543 43772 28552
rect 43720 28509 43729 28543
rect 43729 28509 43763 28543
rect 43763 28509 43772 28543
rect 43720 28500 43772 28509
rect 45008 28543 45060 28552
rect 45008 28509 45017 28543
rect 45017 28509 45051 28543
rect 45051 28509 45060 28543
rect 45008 28500 45060 28509
rect 45836 28568 45888 28620
rect 45560 28500 45612 28552
rect 47952 28568 48004 28620
rect 57796 28611 57848 28620
rect 40224 28432 40276 28484
rect 40684 28475 40736 28484
rect 40684 28441 40693 28475
rect 40693 28441 40727 28475
rect 40727 28441 40736 28475
rect 40684 28432 40736 28441
rect 40776 28432 40828 28484
rect 45284 28475 45336 28484
rect 33140 28364 33192 28416
rect 33508 28407 33560 28416
rect 33508 28373 33517 28407
rect 33517 28373 33551 28407
rect 33551 28373 33560 28407
rect 33508 28364 33560 28373
rect 36176 28364 36228 28416
rect 38108 28364 38160 28416
rect 43904 28407 43956 28416
rect 43904 28373 43913 28407
rect 43913 28373 43947 28407
rect 43947 28373 43956 28407
rect 43904 28364 43956 28373
rect 45284 28441 45293 28475
rect 45293 28441 45327 28475
rect 45327 28441 45336 28475
rect 45284 28432 45336 28441
rect 45376 28475 45428 28484
rect 45376 28441 45393 28475
rect 45393 28441 45427 28475
rect 45427 28441 45428 28475
rect 45376 28432 45428 28441
rect 46020 28432 46072 28484
rect 47216 28500 47268 28552
rect 47768 28543 47820 28552
rect 47768 28509 47777 28543
rect 47777 28509 47811 28543
rect 47811 28509 47820 28543
rect 47768 28500 47820 28509
rect 47860 28543 47912 28552
rect 47860 28509 47869 28543
rect 47869 28509 47903 28543
rect 47903 28509 47912 28543
rect 47860 28500 47912 28509
rect 50160 28543 50212 28552
rect 50160 28509 50169 28543
rect 50169 28509 50203 28543
rect 50203 28509 50212 28543
rect 50160 28500 50212 28509
rect 50620 28500 50672 28552
rect 51908 28500 51960 28552
rect 52460 28543 52512 28552
rect 52460 28509 52466 28543
rect 52466 28509 52500 28543
rect 52500 28509 52512 28543
rect 52460 28500 52512 28509
rect 52920 28543 52972 28552
rect 52920 28509 52929 28543
rect 52929 28509 52963 28543
rect 52963 28509 52972 28543
rect 57796 28577 57805 28611
rect 57805 28577 57839 28611
rect 57839 28577 57848 28611
rect 57796 28568 57848 28577
rect 52920 28500 52972 28509
rect 54668 28500 54720 28552
rect 56324 28543 56376 28552
rect 56324 28509 56333 28543
rect 56333 28509 56367 28543
rect 56367 28509 56376 28543
rect 56324 28500 56376 28509
rect 51632 28475 51684 28484
rect 51632 28441 51641 28475
rect 51641 28441 51675 28475
rect 51675 28441 51684 28475
rect 51632 28432 51684 28441
rect 45192 28364 45244 28416
rect 45652 28407 45704 28416
rect 45652 28373 45661 28407
rect 45661 28373 45695 28407
rect 45695 28373 45704 28407
rect 45652 28364 45704 28373
rect 45836 28364 45888 28416
rect 47584 28364 47636 28416
rect 53196 28432 53248 28484
rect 52368 28364 52420 28416
rect 54392 28432 54444 28484
rect 56968 28432 57020 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 31024 28160 31076 28212
rect 31576 28160 31628 28212
rect 28816 28024 28868 28076
rect 29276 28024 29328 28076
rect 32680 28160 32732 28212
rect 38292 28160 38344 28212
rect 39212 28160 39264 28212
rect 43352 28203 43404 28212
rect 43352 28169 43361 28203
rect 43361 28169 43395 28203
rect 43395 28169 43404 28203
rect 43352 28160 43404 28169
rect 44364 28203 44416 28212
rect 44364 28169 44373 28203
rect 44373 28169 44407 28203
rect 44407 28169 44416 28203
rect 44364 28160 44416 28169
rect 45100 28160 45152 28212
rect 45560 28160 45612 28212
rect 46112 28160 46164 28212
rect 47952 28203 48004 28212
rect 47952 28169 47961 28203
rect 47961 28169 47995 28203
rect 47995 28169 48004 28203
rect 47952 28160 48004 28169
rect 48320 28160 48372 28212
rect 49608 28203 49660 28212
rect 49608 28169 49617 28203
rect 49617 28169 49651 28203
rect 49651 28169 49660 28203
rect 49608 28160 49660 28169
rect 50068 28160 50120 28212
rect 53012 28160 53064 28212
rect 31208 28067 31260 28076
rect 29000 27956 29052 28008
rect 29644 27999 29696 28008
rect 29644 27965 29653 27999
rect 29653 27965 29687 27999
rect 29687 27965 29696 27999
rect 29644 27956 29696 27965
rect 31208 28033 31217 28067
rect 31217 28033 31251 28067
rect 31251 28033 31260 28067
rect 31208 28024 31260 28033
rect 31116 27956 31168 28008
rect 31484 28024 31536 28076
rect 31576 28067 31628 28076
rect 31576 28033 31585 28067
rect 31585 28033 31619 28067
rect 31619 28033 31628 28067
rect 31576 28024 31628 28033
rect 33048 28067 33100 28076
rect 33048 28033 33057 28067
rect 33057 28033 33091 28067
rect 33091 28033 33100 28067
rect 33048 28024 33100 28033
rect 32220 27999 32272 28008
rect 32220 27965 32229 27999
rect 32229 27965 32263 27999
rect 32263 27965 32272 27999
rect 32220 27956 32272 27965
rect 32680 27956 32732 28008
rect 33508 28092 33560 28144
rect 34060 28135 34112 28144
rect 34060 28101 34094 28135
rect 34094 28101 34112 28135
rect 34060 28092 34112 28101
rect 33784 28067 33836 28076
rect 33784 28033 33793 28067
rect 33793 28033 33827 28067
rect 33827 28033 33836 28067
rect 33784 28024 33836 28033
rect 36176 28024 36228 28076
rect 36360 28067 36412 28076
rect 36360 28033 36369 28067
rect 36369 28033 36403 28067
rect 36403 28033 36412 28067
rect 36360 28024 36412 28033
rect 37740 28092 37792 28144
rect 37280 28067 37332 28076
rect 37280 28033 37289 28067
rect 37289 28033 37323 28067
rect 37323 28033 37332 28067
rect 37280 28024 37332 28033
rect 37464 28024 37516 28076
rect 37924 28024 37976 28076
rect 38384 28024 38436 28076
rect 39212 28067 39264 28076
rect 39212 28033 39221 28067
rect 39221 28033 39255 28067
rect 39255 28033 39264 28067
rect 39212 28024 39264 28033
rect 40960 28092 41012 28144
rect 43444 28092 43496 28144
rect 45376 28092 45428 28144
rect 47216 28092 47268 28144
rect 29368 27888 29420 27940
rect 29828 27888 29880 27940
rect 29000 27820 29052 27872
rect 29276 27820 29328 27872
rect 37188 27888 37240 27940
rect 39028 27888 39080 27940
rect 32128 27863 32180 27872
rect 32128 27829 32137 27863
rect 32137 27829 32171 27863
rect 32171 27829 32180 27863
rect 32128 27820 32180 27829
rect 34428 27820 34480 27872
rect 36544 27820 36596 27872
rect 37740 27820 37792 27872
rect 37832 27820 37884 27872
rect 43260 28024 43312 28076
rect 44732 28024 44784 28076
rect 43904 27999 43956 28008
rect 43904 27965 43913 27999
rect 43913 27965 43947 27999
rect 43947 27965 43956 27999
rect 43904 27956 43956 27965
rect 46388 28024 46440 28076
rect 46480 28067 46532 28076
rect 46480 28033 46489 28067
rect 46489 28033 46523 28067
rect 46523 28033 46532 28067
rect 46480 28024 46532 28033
rect 46664 28067 46716 28076
rect 46664 28033 46673 28067
rect 46673 28033 46707 28067
rect 46707 28033 46716 28067
rect 47860 28092 47912 28144
rect 53472 28160 53524 28212
rect 55496 28160 55548 28212
rect 46664 28024 46716 28033
rect 48044 28024 48096 28076
rect 48872 28024 48924 28076
rect 45836 27956 45888 28008
rect 47492 27956 47544 28008
rect 45192 27888 45244 27940
rect 48964 27888 49016 27940
rect 49884 28024 49936 28076
rect 50068 27999 50120 28008
rect 50068 27965 50077 27999
rect 50077 27965 50111 27999
rect 50111 27965 50120 27999
rect 50068 27956 50120 27965
rect 49608 27888 49660 27940
rect 51080 28024 51132 28076
rect 51632 28067 51684 28076
rect 51632 28033 51641 28067
rect 51641 28033 51675 28067
rect 51675 28033 51684 28067
rect 51632 28024 51684 28033
rect 51356 27956 51408 28008
rect 52828 28024 52880 28076
rect 54484 28067 54536 28076
rect 52368 27956 52420 28008
rect 53104 27999 53156 28008
rect 53104 27965 53113 27999
rect 53113 27965 53147 27999
rect 53147 27965 53156 27999
rect 53104 27956 53156 27965
rect 51908 27888 51960 27940
rect 54484 28033 54493 28067
rect 54493 28033 54527 28067
rect 54527 28033 54536 28067
rect 54484 28024 54536 28033
rect 54668 28067 54720 28076
rect 54668 28033 54677 28067
rect 54677 28033 54711 28067
rect 54711 28033 54720 28067
rect 54668 28024 54720 28033
rect 56324 28024 56376 28076
rect 43812 27820 43864 27872
rect 43904 27820 43956 27872
rect 45284 27820 45336 27872
rect 47768 27863 47820 27872
rect 47768 27829 47777 27863
rect 47777 27829 47811 27863
rect 47811 27829 47820 27863
rect 47768 27820 47820 27829
rect 52460 27820 52512 27872
rect 53104 27820 53156 27872
rect 53656 27820 53708 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 28816 27659 28868 27668
rect 28816 27625 28825 27659
rect 28825 27625 28859 27659
rect 28859 27625 28868 27659
rect 28816 27616 28868 27625
rect 31668 27616 31720 27668
rect 31852 27616 31904 27668
rect 31576 27548 31628 27600
rect 31760 27548 31812 27600
rect 1952 27412 2004 27464
rect 29276 27480 29328 27532
rect 29092 27412 29144 27464
rect 28724 27344 28776 27396
rect 31300 27480 31352 27532
rect 32036 27480 32088 27532
rect 30472 27455 30524 27464
rect 30472 27421 30481 27455
rect 30481 27421 30515 27455
rect 30515 27421 30524 27455
rect 30472 27412 30524 27421
rect 30748 27412 30800 27464
rect 29828 27387 29880 27396
rect 29828 27353 29837 27387
rect 29837 27353 29871 27387
rect 29871 27353 29880 27387
rect 29828 27344 29880 27353
rect 30288 27344 30340 27396
rect 31484 27412 31536 27464
rect 31576 27412 31628 27464
rect 33048 27616 33100 27668
rect 36360 27616 36412 27668
rect 37188 27616 37240 27668
rect 38016 27616 38068 27668
rect 38200 27616 38252 27668
rect 41052 27616 41104 27668
rect 41696 27616 41748 27668
rect 43720 27616 43772 27668
rect 32864 27548 32916 27600
rect 36176 27548 36228 27600
rect 38016 27480 38068 27532
rect 44732 27548 44784 27600
rect 45192 27616 45244 27668
rect 45928 27616 45980 27668
rect 46388 27659 46440 27668
rect 46388 27625 46397 27659
rect 46397 27625 46431 27659
rect 46431 27625 46440 27659
rect 46388 27616 46440 27625
rect 47768 27616 47820 27668
rect 47860 27616 47912 27668
rect 52920 27659 52972 27668
rect 52920 27625 52929 27659
rect 52929 27625 52963 27659
rect 52963 27625 52972 27659
rect 52920 27616 52972 27625
rect 48872 27548 48924 27600
rect 31944 27344 31996 27396
rect 36360 27455 36412 27464
rect 32496 27387 32548 27396
rect 32496 27353 32505 27387
rect 32505 27353 32539 27387
rect 32539 27353 32548 27387
rect 36360 27421 36369 27455
rect 36369 27421 36403 27455
rect 36403 27421 36412 27455
rect 36360 27412 36412 27421
rect 37096 27455 37148 27464
rect 37096 27421 37105 27455
rect 37105 27421 37139 27455
rect 37139 27421 37148 27455
rect 37096 27412 37148 27421
rect 37372 27412 37424 27464
rect 37648 27412 37700 27464
rect 37832 27412 37884 27464
rect 41512 27455 41564 27464
rect 41512 27421 41521 27455
rect 41521 27421 41555 27455
rect 41555 27421 41564 27455
rect 41788 27455 41840 27464
rect 41512 27412 41564 27421
rect 41788 27421 41797 27455
rect 41797 27421 41831 27455
rect 41831 27421 41840 27455
rect 41788 27412 41840 27421
rect 42340 27455 42392 27464
rect 42340 27421 42349 27455
rect 42349 27421 42383 27455
rect 42383 27421 42392 27455
rect 42340 27412 42392 27421
rect 43904 27412 43956 27464
rect 45192 27455 45244 27464
rect 45192 27421 45201 27455
rect 45201 27421 45235 27455
rect 45235 27421 45244 27455
rect 45192 27412 45244 27421
rect 45744 27412 45796 27464
rect 45928 27455 45980 27464
rect 45928 27421 45937 27455
rect 45937 27421 45971 27455
rect 45971 27421 45980 27455
rect 45928 27412 45980 27421
rect 32496 27344 32548 27353
rect 30380 27276 30432 27328
rect 32128 27276 32180 27328
rect 32864 27319 32916 27328
rect 32864 27285 32873 27319
rect 32873 27285 32907 27319
rect 32907 27285 32916 27319
rect 32864 27276 32916 27285
rect 36728 27276 36780 27328
rect 38292 27344 38344 27396
rect 41696 27387 41748 27396
rect 41696 27353 41705 27387
rect 41705 27353 41739 27387
rect 41739 27353 41748 27387
rect 41696 27344 41748 27353
rect 42800 27344 42852 27396
rect 43260 27344 43312 27396
rect 39488 27276 39540 27328
rect 40592 27276 40644 27328
rect 42340 27276 42392 27328
rect 45376 27319 45428 27328
rect 45376 27285 45385 27319
rect 45385 27285 45419 27319
rect 45419 27285 45428 27319
rect 45376 27276 45428 27285
rect 45928 27276 45980 27328
rect 47676 27480 47728 27532
rect 56968 27591 57020 27600
rect 46296 27412 46348 27464
rect 47308 27455 47360 27464
rect 47308 27421 47317 27455
rect 47317 27421 47351 27455
rect 47351 27421 47360 27455
rect 48136 27455 48188 27464
rect 47308 27412 47360 27421
rect 48136 27421 48145 27455
rect 48145 27421 48179 27455
rect 48179 27421 48188 27455
rect 48136 27412 48188 27421
rect 48320 27412 48372 27464
rect 49424 27455 49476 27464
rect 49424 27421 49433 27455
rect 49433 27421 49467 27455
rect 49467 27421 49476 27455
rect 49884 27480 49936 27532
rect 56968 27557 56977 27591
rect 56977 27557 57011 27591
rect 57011 27557 57020 27591
rect 56968 27548 57020 27557
rect 49424 27412 49476 27421
rect 51448 27455 51500 27464
rect 51448 27421 51457 27455
rect 51457 27421 51491 27455
rect 51491 27421 51500 27455
rect 51448 27412 51500 27421
rect 49240 27387 49292 27396
rect 49240 27353 49249 27387
rect 49249 27353 49283 27387
rect 49283 27353 49292 27387
rect 49240 27344 49292 27353
rect 49608 27344 49660 27396
rect 50804 27344 50856 27396
rect 50160 27276 50212 27328
rect 51172 27344 51224 27396
rect 52368 27412 52420 27464
rect 53012 27480 53064 27532
rect 54484 27480 54536 27532
rect 53196 27412 53248 27464
rect 53656 27455 53708 27464
rect 53656 27421 53665 27455
rect 53665 27421 53699 27455
rect 53699 27421 53708 27455
rect 53656 27412 53708 27421
rect 56784 27412 56836 27464
rect 51540 27276 51592 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 8484 27072 8536 27124
rect 29828 27072 29880 27124
rect 30748 27072 30800 27124
rect 31484 27072 31536 27124
rect 37740 27115 37792 27124
rect 37740 27081 37749 27115
rect 37749 27081 37783 27115
rect 37783 27081 37792 27115
rect 37740 27072 37792 27081
rect 30472 27004 30524 27056
rect 1952 26979 2004 26988
rect 1952 26945 1961 26979
rect 1961 26945 1995 26979
rect 1995 26945 2004 26979
rect 1952 26936 2004 26945
rect 8760 26979 8812 26988
rect 8760 26945 8769 26979
rect 8769 26945 8803 26979
rect 8803 26945 8812 26979
rect 8760 26936 8812 26945
rect 2504 26868 2556 26920
rect 2780 26911 2832 26920
rect 2780 26877 2789 26911
rect 2789 26877 2823 26911
rect 2823 26877 2832 26911
rect 2780 26868 2832 26877
rect 8576 26868 8628 26920
rect 29000 26868 29052 26920
rect 28816 26800 28868 26852
rect 29552 26936 29604 26988
rect 29736 26936 29788 26988
rect 31300 27004 31352 27056
rect 32128 27047 32180 27056
rect 31116 26936 31168 26988
rect 32128 27013 32137 27047
rect 32137 27013 32171 27047
rect 32171 27013 32180 27047
rect 32128 27004 32180 27013
rect 36820 27004 36872 27056
rect 36728 26979 36780 26988
rect 36728 26945 36737 26979
rect 36737 26945 36771 26979
rect 36771 26945 36780 26979
rect 36728 26936 36780 26945
rect 38844 27004 38896 27056
rect 37832 26979 37884 26988
rect 37832 26945 37841 26979
rect 37841 26945 37875 26979
rect 37875 26945 37884 26979
rect 37832 26936 37884 26945
rect 38384 26936 38436 26988
rect 40500 27004 40552 27056
rect 29644 26868 29696 26920
rect 30012 26868 30064 26920
rect 30932 26868 30984 26920
rect 31208 26911 31260 26920
rect 31208 26877 31217 26911
rect 31217 26877 31251 26911
rect 31251 26877 31260 26911
rect 31208 26868 31260 26877
rect 31300 26868 31352 26920
rect 32496 26868 32548 26920
rect 37648 26868 37700 26920
rect 30840 26800 30892 26852
rect 32220 26800 32272 26852
rect 36544 26800 36596 26852
rect 40684 26936 40736 26988
rect 41052 26936 41104 26988
rect 41512 27072 41564 27124
rect 44640 27072 44692 27124
rect 48136 27072 48188 27124
rect 49332 27072 49384 27124
rect 51356 27072 51408 27124
rect 51540 27115 51592 27124
rect 51540 27081 51549 27115
rect 51549 27081 51583 27115
rect 51583 27081 51592 27115
rect 51540 27072 51592 27081
rect 51908 27072 51960 27124
rect 55956 27072 56008 27124
rect 41236 27047 41288 27056
rect 41236 27013 41245 27047
rect 41245 27013 41279 27047
rect 41279 27013 41288 27047
rect 41236 27004 41288 27013
rect 42340 27004 42392 27056
rect 42800 26936 42852 26988
rect 43720 26979 43772 26988
rect 43720 26945 43729 26979
rect 43729 26945 43763 26979
rect 43763 26945 43772 26979
rect 43720 26936 43772 26945
rect 46296 26979 46348 26988
rect 40224 26868 40276 26920
rect 43536 26868 43588 26920
rect 46296 26945 46305 26979
rect 46305 26945 46339 26979
rect 46339 26945 46348 26979
rect 46296 26936 46348 26945
rect 47308 27004 47360 27056
rect 48964 27004 49016 27056
rect 49884 27004 49936 27056
rect 51632 27004 51684 27056
rect 48044 26979 48096 26988
rect 48044 26945 48053 26979
rect 48053 26945 48087 26979
rect 48087 26945 48096 26979
rect 48044 26936 48096 26945
rect 47124 26868 47176 26920
rect 56600 26936 56652 26988
rect 49700 26911 49752 26920
rect 49700 26877 49709 26911
rect 49709 26877 49743 26911
rect 49743 26877 49752 26911
rect 49700 26868 49752 26877
rect 50344 26868 50396 26920
rect 50712 26868 50764 26920
rect 51448 26868 51500 26920
rect 40040 26800 40092 26852
rect 49240 26800 49292 26852
rect 50160 26800 50212 26852
rect 51080 26843 51132 26852
rect 51080 26809 51089 26843
rect 51089 26809 51123 26843
rect 51123 26809 51132 26843
rect 51080 26800 51132 26809
rect 30656 26732 30708 26784
rect 38752 26732 38804 26784
rect 40408 26732 40460 26784
rect 44088 26732 44140 26784
rect 47676 26732 47728 26784
rect 49332 26732 49384 26784
rect 50344 26732 50396 26784
rect 52460 26732 52512 26784
rect 56968 26732 57020 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2504 26571 2556 26580
rect 2504 26537 2513 26571
rect 2513 26537 2547 26571
rect 2547 26537 2556 26571
rect 2504 26528 2556 26537
rect 47124 26528 47176 26580
rect 47216 26528 47268 26580
rect 50160 26528 50212 26580
rect 51632 26528 51684 26580
rect 8760 26324 8812 26376
rect 9220 26324 9272 26376
rect 20260 26324 20312 26376
rect 24860 26324 24912 26376
rect 29368 26324 29420 26376
rect 29736 26367 29788 26376
rect 29736 26333 29745 26367
rect 29745 26333 29779 26367
rect 29779 26333 29788 26367
rect 29736 26324 29788 26333
rect 30012 26324 30064 26376
rect 30288 26324 30340 26376
rect 30840 26392 30892 26444
rect 32036 26460 32088 26512
rect 32128 26460 32180 26512
rect 37096 26460 37148 26512
rect 30748 26367 30800 26376
rect 30748 26333 30757 26367
rect 30757 26333 30791 26367
rect 30791 26333 30800 26367
rect 30748 26324 30800 26333
rect 30932 26367 30984 26376
rect 30932 26333 30941 26367
rect 30941 26333 30975 26367
rect 30975 26333 30984 26367
rect 30932 26324 30984 26333
rect 28816 26256 28868 26308
rect 30196 26256 30248 26308
rect 31668 26324 31720 26376
rect 31300 26256 31352 26308
rect 31208 26188 31260 26240
rect 31852 26367 31904 26376
rect 31852 26333 31861 26367
rect 31861 26333 31895 26367
rect 31895 26333 31904 26367
rect 31852 26324 31904 26333
rect 31944 26256 31996 26308
rect 32220 26324 32272 26376
rect 39212 26460 39264 26512
rect 40316 26460 40368 26512
rect 38752 26392 38804 26444
rect 43444 26460 43496 26512
rect 44456 26460 44508 26512
rect 37832 26367 37884 26376
rect 37832 26333 37841 26367
rect 37841 26333 37875 26367
rect 37875 26333 37884 26367
rect 37832 26324 37884 26333
rect 40040 26367 40092 26376
rect 40040 26333 40049 26367
rect 40049 26333 40083 26367
rect 40083 26333 40092 26367
rect 40040 26324 40092 26333
rect 43720 26392 43772 26444
rect 40592 26324 40644 26376
rect 41420 26367 41472 26376
rect 41420 26333 41429 26367
rect 41429 26333 41463 26367
rect 41463 26333 41472 26367
rect 41420 26324 41472 26333
rect 41604 26367 41656 26376
rect 41604 26333 41613 26367
rect 41613 26333 41647 26367
rect 41647 26333 41656 26367
rect 41604 26324 41656 26333
rect 41788 26324 41840 26376
rect 43076 26367 43128 26376
rect 43076 26333 43085 26367
rect 43085 26333 43119 26367
rect 43119 26333 43128 26367
rect 43076 26324 43128 26333
rect 44180 26324 44232 26376
rect 38660 26256 38712 26308
rect 38844 26256 38896 26308
rect 40500 26256 40552 26308
rect 37280 26188 37332 26240
rect 38108 26188 38160 26240
rect 39764 26188 39816 26240
rect 41880 26256 41932 26308
rect 43812 26256 43864 26308
rect 41696 26188 41748 26240
rect 42800 26188 42852 26240
rect 43996 26188 44048 26240
rect 44640 26256 44692 26308
rect 50712 26460 50764 26512
rect 51080 26392 51132 26444
rect 56968 26392 57020 26444
rect 58164 26435 58216 26444
rect 58164 26401 58173 26435
rect 58173 26401 58207 26435
rect 58207 26401 58216 26435
rect 58164 26392 58216 26401
rect 48964 26324 49016 26376
rect 50160 26367 50212 26376
rect 50160 26333 50169 26367
rect 50169 26333 50203 26367
rect 50203 26333 50212 26367
rect 50160 26324 50212 26333
rect 50344 26367 50396 26376
rect 50344 26333 50353 26367
rect 50353 26333 50387 26367
rect 50387 26333 50396 26367
rect 50344 26324 50396 26333
rect 50620 26324 50672 26376
rect 46388 26256 46440 26308
rect 49884 26256 49936 26308
rect 51264 26299 51316 26308
rect 51264 26265 51305 26299
rect 51305 26265 51316 26299
rect 51264 26256 51316 26265
rect 52276 26256 52328 26308
rect 57060 26256 57112 26308
rect 47676 26188 47728 26240
rect 48044 26188 48096 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 37372 25984 37424 26036
rect 40868 25984 40920 26036
rect 43720 25984 43772 26036
rect 46296 25984 46348 26036
rect 49240 25984 49292 26036
rect 51264 25984 51316 26036
rect 57060 26027 57112 26036
rect 57060 25993 57069 26027
rect 57069 25993 57103 26027
rect 57103 25993 57112 26027
rect 57060 25984 57112 25993
rect 2688 25916 2740 25968
rect 9864 25916 9916 25968
rect 16580 25916 16632 25968
rect 39580 25916 39632 25968
rect 8760 25891 8812 25900
rect 8760 25857 8769 25891
rect 8769 25857 8803 25891
rect 8803 25857 8812 25891
rect 8760 25848 8812 25857
rect 30380 25891 30432 25900
rect 30380 25857 30389 25891
rect 30389 25857 30423 25891
rect 30423 25857 30432 25891
rect 30380 25848 30432 25857
rect 30656 25891 30708 25900
rect 9496 25780 9548 25832
rect 26976 25780 27028 25832
rect 29552 25780 29604 25832
rect 30656 25857 30665 25891
rect 30665 25857 30699 25891
rect 30699 25857 30708 25891
rect 30656 25848 30708 25857
rect 31208 25891 31260 25900
rect 31208 25857 31217 25891
rect 31217 25857 31251 25891
rect 31251 25857 31260 25891
rect 31208 25848 31260 25857
rect 31484 25848 31536 25900
rect 37280 25891 37332 25900
rect 37280 25857 37289 25891
rect 37289 25857 37323 25891
rect 37323 25857 37332 25891
rect 37280 25848 37332 25857
rect 37556 25891 37608 25900
rect 37556 25857 37565 25891
rect 37565 25857 37599 25891
rect 37599 25857 37608 25891
rect 37556 25848 37608 25857
rect 37648 25848 37700 25900
rect 38016 25891 38068 25900
rect 38016 25857 38025 25891
rect 38025 25857 38059 25891
rect 38059 25857 38068 25891
rect 38016 25848 38068 25857
rect 38936 25891 38988 25900
rect 38936 25857 38945 25891
rect 38945 25857 38979 25891
rect 38979 25857 38988 25891
rect 38936 25848 38988 25857
rect 39488 25848 39540 25900
rect 39856 25925 39908 25934
rect 39856 25891 39865 25925
rect 39865 25891 39899 25925
rect 39899 25891 39908 25925
rect 40316 25916 40368 25968
rect 39856 25882 39908 25891
rect 40040 25848 40092 25900
rect 32864 25780 32916 25832
rect 38752 25823 38804 25832
rect 38752 25789 38761 25823
rect 38761 25789 38795 25823
rect 38795 25789 38804 25823
rect 38752 25780 38804 25789
rect 38844 25823 38896 25832
rect 38844 25789 38853 25823
rect 38853 25789 38887 25823
rect 38887 25789 38896 25823
rect 38844 25780 38896 25789
rect 40592 25848 40644 25900
rect 40868 25848 40920 25900
rect 41604 25891 41656 25900
rect 41604 25857 41613 25891
rect 41613 25857 41647 25891
rect 41647 25857 41656 25891
rect 41604 25848 41656 25857
rect 41788 25891 41840 25900
rect 41788 25857 41797 25891
rect 41797 25857 41831 25891
rect 41831 25857 41840 25891
rect 41788 25848 41840 25857
rect 43444 25891 43496 25900
rect 29368 25644 29420 25696
rect 31024 25644 31076 25696
rect 38292 25644 38344 25696
rect 40316 25780 40368 25832
rect 41420 25780 41472 25832
rect 43444 25857 43453 25891
rect 43453 25857 43487 25891
rect 43487 25857 43496 25891
rect 43444 25848 43496 25857
rect 43536 25848 43588 25900
rect 44364 25848 44416 25900
rect 48872 25891 48924 25900
rect 48872 25857 48881 25891
rect 48881 25857 48915 25891
rect 48915 25857 48924 25891
rect 48872 25848 48924 25857
rect 44272 25823 44324 25832
rect 44272 25789 44281 25823
rect 44281 25789 44315 25823
rect 44315 25789 44324 25823
rect 44272 25780 44324 25789
rect 44088 25712 44140 25764
rect 49700 25848 49752 25900
rect 57428 25848 57480 25900
rect 40408 25644 40460 25696
rect 40684 25644 40736 25696
rect 41696 25644 41748 25696
rect 47768 25644 47820 25696
rect 49240 25687 49292 25696
rect 49240 25653 49249 25687
rect 49249 25653 49283 25687
rect 49283 25653 49292 25687
rect 49240 25644 49292 25653
rect 56508 25644 56560 25696
rect 58072 25687 58124 25696
rect 58072 25653 58081 25687
rect 58081 25653 58115 25687
rect 58115 25653 58124 25687
rect 58072 25644 58124 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 40040 25440 40092 25492
rect 42800 25440 42852 25492
rect 44364 25440 44416 25492
rect 45284 25440 45336 25492
rect 37096 25304 37148 25356
rect 38752 25372 38804 25424
rect 39120 25372 39172 25424
rect 40132 25372 40184 25424
rect 39488 25304 39540 25356
rect 8760 25236 8812 25288
rect 37280 25236 37332 25288
rect 38016 25236 38068 25288
rect 38292 25279 38344 25288
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 9864 25211 9916 25220
rect 9864 25177 9873 25211
rect 9873 25177 9907 25211
rect 9907 25177 9916 25211
rect 9864 25168 9916 25177
rect 38844 25236 38896 25288
rect 39120 25279 39172 25288
rect 39120 25245 39129 25279
rect 39129 25245 39163 25279
rect 39163 25245 39172 25279
rect 39120 25236 39172 25245
rect 39764 25168 39816 25220
rect 40316 25279 40368 25288
rect 40316 25245 40325 25279
rect 40325 25245 40359 25279
rect 40359 25245 40368 25279
rect 40316 25236 40368 25245
rect 40500 25236 40552 25288
rect 41144 25279 41196 25288
rect 41144 25245 41153 25279
rect 41153 25245 41187 25279
rect 41187 25245 41196 25279
rect 41144 25236 41196 25245
rect 41236 25236 41288 25288
rect 42708 25279 42760 25288
rect 42708 25245 42717 25279
rect 42717 25245 42751 25279
rect 42751 25245 42760 25279
rect 42708 25236 42760 25245
rect 44180 25372 44232 25424
rect 42892 25279 42944 25288
rect 42892 25245 42901 25279
rect 42901 25245 42935 25279
rect 42935 25245 42944 25279
rect 42892 25236 42944 25245
rect 43076 25279 43128 25288
rect 43076 25245 43085 25279
rect 43085 25245 43119 25279
rect 43119 25245 43128 25279
rect 43076 25236 43128 25245
rect 43444 25236 43496 25288
rect 47676 25304 47728 25356
rect 58072 25372 58124 25424
rect 56508 25347 56560 25356
rect 56508 25313 56517 25347
rect 56517 25313 56551 25347
rect 56551 25313 56560 25347
rect 56508 25304 56560 25313
rect 58164 25347 58216 25356
rect 58164 25313 58173 25347
rect 58173 25313 58207 25347
rect 58207 25313 58216 25347
rect 58164 25304 58216 25313
rect 47768 25279 47820 25288
rect 37832 25143 37884 25152
rect 37832 25109 37841 25143
rect 37841 25109 37875 25143
rect 37875 25109 37884 25143
rect 37832 25100 37884 25109
rect 39120 25100 39172 25152
rect 40224 25100 40276 25152
rect 40960 25168 41012 25220
rect 41972 25211 42024 25220
rect 41972 25177 41981 25211
rect 41981 25177 42015 25211
rect 42015 25177 42024 25211
rect 41972 25168 42024 25177
rect 44088 25211 44140 25220
rect 44088 25177 44097 25211
rect 44097 25177 44131 25211
rect 44131 25177 44140 25211
rect 44088 25168 44140 25177
rect 47768 25245 47777 25279
rect 47777 25245 47811 25279
rect 47811 25245 47820 25279
rect 47768 25236 47820 25245
rect 48872 25236 48924 25288
rect 41420 25100 41472 25152
rect 41788 25100 41840 25152
rect 43996 25100 44048 25152
rect 44272 25143 44324 25152
rect 44272 25109 44297 25143
rect 44297 25109 44324 25143
rect 45192 25143 45244 25152
rect 44272 25100 44324 25109
rect 45192 25109 45201 25143
rect 45201 25109 45235 25143
rect 45235 25109 45244 25143
rect 45192 25100 45244 25109
rect 47308 25143 47360 25152
rect 47308 25109 47317 25143
rect 47317 25109 47351 25143
rect 47351 25109 47360 25143
rect 47308 25100 47360 25109
rect 47676 25100 47728 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 38660 24939 38712 24948
rect 38660 24905 38669 24939
rect 38669 24905 38703 24939
rect 38703 24905 38712 24939
rect 38660 24896 38712 24905
rect 38844 24896 38896 24948
rect 41420 24896 41472 24948
rect 37832 24828 37884 24880
rect 2320 24803 2372 24812
rect 2320 24769 2329 24803
rect 2329 24769 2363 24803
rect 2363 24769 2372 24803
rect 2320 24760 2372 24769
rect 8576 24760 8628 24812
rect 8760 24803 8812 24812
rect 8760 24769 8769 24803
rect 8769 24769 8803 24803
rect 8803 24769 8812 24803
rect 8760 24760 8812 24769
rect 37556 24803 37608 24812
rect 37556 24769 37565 24803
rect 37565 24769 37599 24803
rect 37599 24769 37608 24803
rect 37556 24760 37608 24769
rect 38108 24760 38160 24812
rect 40500 24828 40552 24880
rect 41236 24871 41288 24880
rect 41236 24837 41245 24871
rect 41245 24837 41279 24871
rect 41279 24837 41288 24871
rect 41236 24828 41288 24837
rect 9036 24735 9088 24744
rect 9036 24701 9045 24735
rect 9045 24701 9079 24735
rect 9079 24701 9088 24735
rect 9036 24692 9088 24701
rect 38844 24760 38896 24812
rect 39120 24760 39172 24812
rect 41052 24803 41104 24812
rect 41052 24769 41061 24803
rect 41061 24769 41095 24803
rect 41095 24769 41104 24803
rect 41052 24760 41104 24769
rect 40316 24735 40368 24744
rect 40316 24701 40325 24735
rect 40325 24701 40359 24735
rect 40359 24701 40368 24735
rect 40316 24692 40368 24701
rect 38660 24624 38712 24676
rect 1952 24556 2004 24608
rect 2136 24556 2188 24608
rect 39304 24556 39356 24608
rect 40960 24624 41012 24676
rect 41420 24803 41472 24812
rect 41420 24769 41429 24803
rect 41429 24769 41463 24803
rect 41463 24769 41472 24803
rect 41420 24760 41472 24769
rect 42892 24896 42944 24948
rect 45192 24896 45244 24948
rect 47216 24896 47268 24948
rect 44640 24828 44692 24880
rect 46296 24828 46348 24880
rect 42984 24760 43036 24812
rect 41880 24692 41932 24744
rect 44548 24735 44600 24744
rect 44548 24701 44557 24735
rect 44557 24701 44591 24735
rect 44591 24701 44600 24735
rect 44548 24692 44600 24701
rect 45284 24803 45336 24812
rect 45284 24769 45293 24803
rect 45293 24769 45327 24803
rect 45327 24769 45336 24803
rect 45284 24760 45336 24769
rect 46388 24760 46440 24812
rect 42800 24667 42852 24676
rect 40132 24556 40184 24608
rect 42800 24633 42809 24667
rect 42809 24633 42843 24667
rect 42843 24633 42852 24667
rect 42800 24624 42852 24633
rect 43628 24667 43680 24676
rect 43628 24633 43637 24667
rect 43637 24633 43671 24667
rect 43671 24633 43680 24667
rect 43628 24624 43680 24633
rect 43996 24624 44048 24676
rect 44732 24624 44784 24676
rect 43444 24556 43496 24608
rect 44916 24556 44968 24608
rect 45468 24624 45520 24676
rect 46756 24803 46808 24812
rect 46756 24769 46765 24803
rect 46765 24769 46799 24803
rect 46799 24769 46808 24803
rect 46756 24760 46808 24769
rect 47584 24803 47636 24812
rect 47584 24769 47593 24803
rect 47593 24769 47627 24803
rect 47627 24769 47636 24803
rect 47584 24760 47636 24769
rect 56600 24760 56652 24812
rect 57428 24760 57480 24812
rect 46664 24624 46716 24676
rect 47216 24624 47268 24676
rect 45744 24599 45796 24608
rect 45744 24565 45753 24599
rect 45753 24565 45787 24599
rect 45787 24565 45796 24599
rect 45744 24556 45796 24565
rect 45836 24556 45888 24608
rect 47952 24735 48004 24744
rect 47952 24701 47961 24735
rect 47961 24701 47995 24735
rect 47995 24701 48004 24735
rect 47952 24692 48004 24701
rect 47584 24624 47636 24676
rect 49240 24624 49292 24676
rect 47676 24599 47728 24608
rect 47676 24565 47685 24599
rect 47685 24565 47719 24599
rect 47719 24565 47728 24599
rect 47676 24556 47728 24565
rect 56508 24556 56560 24608
rect 58072 24599 58124 24608
rect 58072 24565 58081 24599
rect 58081 24565 58115 24599
rect 58115 24565 58124 24599
rect 58072 24556 58124 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 40316 24395 40368 24404
rect 40316 24361 40325 24395
rect 40325 24361 40359 24395
rect 40359 24361 40368 24395
rect 40316 24352 40368 24361
rect 44548 24352 44600 24404
rect 46480 24352 46532 24404
rect 41972 24284 42024 24336
rect 42800 24284 42852 24336
rect 43076 24284 43128 24336
rect 45836 24284 45888 24336
rect 46940 24284 46992 24336
rect 32036 24216 32088 24268
rect 39304 24148 39356 24200
rect 40224 24216 40276 24268
rect 40132 24191 40184 24200
rect 40132 24157 40141 24191
rect 40141 24157 40175 24191
rect 40175 24157 40184 24191
rect 40132 24148 40184 24157
rect 41696 24148 41748 24200
rect 41880 24191 41932 24200
rect 41880 24157 41889 24191
rect 41889 24157 41923 24191
rect 41923 24157 41932 24191
rect 41880 24148 41932 24157
rect 32588 24080 32640 24132
rect 34152 24123 34204 24132
rect 34152 24089 34161 24123
rect 34161 24089 34195 24123
rect 34195 24089 34204 24123
rect 34152 24080 34204 24089
rect 41236 24080 41288 24132
rect 42800 24191 42852 24200
rect 42800 24157 42809 24191
rect 42809 24157 42843 24191
rect 42843 24157 42852 24191
rect 42984 24191 43036 24200
rect 42800 24148 42852 24157
rect 42984 24157 42993 24191
rect 42993 24157 43027 24191
rect 43027 24157 43036 24191
rect 42984 24148 43036 24157
rect 41052 24012 41104 24064
rect 42892 24080 42944 24132
rect 43628 24080 43680 24132
rect 45744 24216 45796 24268
rect 46296 24216 46348 24268
rect 47952 24259 48004 24268
rect 47952 24225 47961 24259
rect 47961 24225 47995 24259
rect 47995 24225 48004 24259
rect 47952 24216 48004 24225
rect 45192 24148 45244 24200
rect 45928 24191 45980 24200
rect 45928 24157 45937 24191
rect 45937 24157 45971 24191
rect 45971 24157 45980 24191
rect 45928 24148 45980 24157
rect 47308 24148 47360 24200
rect 58072 24284 58124 24336
rect 56508 24259 56560 24268
rect 56508 24225 56517 24259
rect 56517 24225 56551 24259
rect 56551 24225 56560 24259
rect 56508 24216 56560 24225
rect 58164 24259 58216 24268
rect 58164 24225 58173 24259
rect 58173 24225 58207 24259
rect 58207 24225 58216 24259
rect 58164 24216 58216 24225
rect 46572 24080 46624 24132
rect 44364 24012 44416 24064
rect 45468 24012 45520 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 32588 23851 32640 23860
rect 32588 23817 32597 23851
rect 32597 23817 32631 23851
rect 32631 23817 32640 23851
rect 32588 23808 32640 23817
rect 2136 23783 2188 23792
rect 2136 23749 2145 23783
rect 2145 23749 2179 23783
rect 2179 23749 2188 23783
rect 2136 23740 2188 23749
rect 43260 23740 43312 23792
rect 44272 23808 44324 23860
rect 45192 23851 45244 23860
rect 45192 23817 45201 23851
rect 45201 23817 45235 23851
rect 45235 23817 45244 23851
rect 45192 23808 45244 23817
rect 45468 23808 45520 23860
rect 47952 23851 48004 23860
rect 1952 23715 2004 23724
rect 1952 23681 1961 23715
rect 1961 23681 1995 23715
rect 1995 23681 2004 23715
rect 1952 23672 2004 23681
rect 33140 23672 33192 23724
rect 43352 23715 43404 23724
rect 43352 23681 43361 23715
rect 43361 23681 43395 23715
rect 43395 23681 43404 23715
rect 43352 23672 43404 23681
rect 43812 23672 43864 23724
rect 2780 23647 2832 23656
rect 2780 23613 2789 23647
rect 2789 23613 2823 23647
rect 2823 23613 2832 23647
rect 2780 23604 2832 23613
rect 44364 23715 44416 23724
rect 44364 23681 44373 23715
rect 44373 23681 44407 23715
rect 44407 23681 44416 23715
rect 44640 23715 44692 23724
rect 44364 23672 44416 23681
rect 44640 23681 44649 23715
rect 44649 23681 44683 23715
rect 44683 23681 44692 23715
rect 44640 23672 44692 23681
rect 44732 23715 44784 23724
rect 44732 23681 44741 23715
rect 44741 23681 44775 23715
rect 44775 23681 44784 23715
rect 45468 23715 45520 23724
rect 44732 23672 44784 23681
rect 45468 23681 45477 23715
rect 45477 23681 45511 23715
rect 45511 23681 45520 23715
rect 45468 23672 45520 23681
rect 46388 23740 46440 23792
rect 45928 23672 45980 23724
rect 46664 23715 46716 23724
rect 46664 23681 46673 23715
rect 46673 23681 46707 23715
rect 46707 23681 46716 23715
rect 46664 23672 46716 23681
rect 47124 23740 47176 23792
rect 47308 23672 47360 23724
rect 47952 23817 47961 23851
rect 47961 23817 47995 23851
rect 47995 23817 48004 23851
rect 47952 23808 48004 23817
rect 47768 23715 47820 23724
rect 47768 23681 47777 23715
rect 47777 23681 47811 23715
rect 47811 23681 47820 23715
rect 47768 23672 47820 23681
rect 44272 23536 44324 23588
rect 45652 23647 45704 23656
rect 45652 23613 45661 23647
rect 45661 23613 45695 23647
rect 45695 23613 45704 23647
rect 46572 23647 46624 23656
rect 45652 23604 45704 23613
rect 46572 23613 46581 23647
rect 46581 23613 46615 23647
rect 46615 23613 46624 23647
rect 46572 23604 46624 23613
rect 44640 23468 44692 23520
rect 45652 23468 45704 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 43904 23264 43956 23316
rect 47768 23264 47820 23316
rect 40040 23196 40092 23248
rect 43260 23128 43312 23180
rect 44364 23128 44416 23180
rect 46296 23128 46348 23180
rect 40408 23060 40460 23112
rect 42892 23060 42944 23112
rect 43076 23103 43128 23112
rect 43076 23069 43085 23103
rect 43085 23069 43119 23103
rect 43119 23069 43128 23103
rect 44272 23103 44324 23112
rect 43076 23060 43128 23069
rect 44272 23069 44281 23103
rect 44281 23069 44315 23103
rect 44315 23069 44324 23103
rect 44272 23060 44324 23069
rect 46940 23103 46992 23112
rect 46940 23069 46949 23103
rect 46949 23069 46983 23103
rect 46983 23069 46992 23103
rect 46940 23060 46992 23069
rect 47124 23103 47176 23112
rect 47124 23069 47133 23103
rect 47133 23069 47167 23103
rect 47167 23069 47176 23103
rect 47124 23060 47176 23069
rect 40684 22924 40736 22976
rect 43720 22992 43772 23044
rect 43352 22924 43404 22976
rect 43536 22924 43588 22976
rect 44364 22924 44416 22976
rect 45468 22967 45520 22976
rect 45468 22933 45477 22967
rect 45477 22933 45511 22967
rect 45511 22933 45520 22967
rect 45468 22924 45520 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 43720 22763 43772 22772
rect 43720 22729 43729 22763
rect 43729 22729 43763 22763
rect 43763 22729 43772 22763
rect 43720 22720 43772 22729
rect 45468 22720 45520 22772
rect 43260 22584 43312 22636
rect 43536 22627 43588 22636
rect 43536 22593 43545 22627
rect 43545 22593 43579 22627
rect 43579 22593 43588 22627
rect 43536 22584 43588 22593
rect 44364 22627 44416 22636
rect 44364 22593 44373 22627
rect 44373 22593 44407 22627
rect 44407 22593 44416 22627
rect 44364 22584 44416 22593
rect 45192 22627 45244 22636
rect 45192 22593 45201 22627
rect 45201 22593 45235 22627
rect 45235 22593 45244 22627
rect 45192 22584 45244 22593
rect 57520 22652 57572 22704
rect 44272 22448 44324 22500
rect 57612 22584 57664 22636
rect 56600 22423 56652 22432
rect 56600 22389 56609 22423
rect 56609 22389 56643 22423
rect 56643 22389 56652 22423
rect 56600 22380 56652 22389
rect 57244 22423 57296 22432
rect 57244 22389 57253 22423
rect 57253 22389 57287 22423
rect 57287 22389 57296 22423
rect 57244 22380 57296 22389
rect 57336 22380 57388 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 43260 22176 43312 22228
rect 44640 22176 44692 22228
rect 45192 22176 45244 22228
rect 1952 21972 2004 22024
rect 43812 22040 43864 22092
rect 43536 21947 43588 21956
rect 43536 21913 43566 21947
rect 43566 21913 43588 21947
rect 43536 21904 43588 21913
rect 43812 21904 43864 21956
rect 44272 21836 44324 21888
rect 57336 22108 57388 22160
rect 56600 22040 56652 22092
rect 57888 22083 57940 22092
rect 57888 22049 57897 22083
rect 57897 22049 57931 22083
rect 57931 22049 57940 22083
rect 57888 22040 57940 22049
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 17132 21675 17184 21684
rect 17132 21641 17141 21675
rect 17141 21641 17175 21675
rect 17175 21641 17184 21675
rect 17132 21632 17184 21641
rect 1952 21539 2004 21548
rect 1952 21505 1961 21539
rect 1961 21505 1995 21539
rect 1995 21505 2004 21539
rect 1952 21496 2004 21505
rect 17408 21496 17460 21548
rect 19432 21496 19484 21548
rect 29644 21496 29696 21548
rect 2136 21471 2188 21480
rect 2136 21437 2145 21471
rect 2145 21437 2179 21471
rect 2179 21437 2188 21471
rect 2136 21428 2188 21437
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 2780 21428 2832 21437
rect 20260 21428 20312 21480
rect 57704 21496 57756 21548
rect 3884 21292 3936 21344
rect 57060 21335 57112 21344
rect 57060 21301 57069 21335
rect 57069 21301 57103 21335
rect 57103 21301 57112 21335
rect 57060 21292 57112 21301
rect 57152 21292 57204 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1952 20884 2004 20936
rect 19432 20884 19484 20936
rect 31208 20952 31260 21004
rect 35348 20952 35400 21004
rect 57888 20995 57940 21004
rect 28448 20884 28500 20936
rect 57888 20961 57897 20995
rect 57897 20961 57931 20995
rect 57931 20961 57940 20995
rect 57888 20952 57940 20961
rect 19340 20748 19392 20800
rect 29644 20816 29696 20868
rect 58072 20884 58124 20936
rect 57244 20816 57296 20868
rect 47584 20748 47636 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 30472 20476 30524 20528
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 19432 20408 19484 20460
rect 29644 20451 29696 20460
rect 29644 20417 29653 20451
rect 29653 20417 29687 20451
rect 29687 20417 29696 20451
rect 29644 20408 29696 20417
rect 58072 20451 58124 20460
rect 58072 20417 58081 20451
rect 58081 20417 58115 20451
rect 58115 20417 58124 20451
rect 58072 20408 58124 20417
rect 2504 20340 2556 20392
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 3976 20340 4028 20392
rect 20352 20383 20404 20392
rect 20352 20349 20361 20383
rect 20361 20349 20395 20383
rect 20395 20349 20404 20383
rect 20352 20340 20404 20349
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2136 20000 2188 20052
rect 31116 19907 31168 19916
rect 31116 19873 31125 19907
rect 31125 19873 31159 19907
rect 31159 19873 31168 19907
rect 57152 19932 57204 19984
rect 31116 19864 31168 19873
rect 2688 19796 2740 19848
rect 19340 19796 19392 19848
rect 19432 19796 19484 19848
rect 29644 19796 29696 19848
rect 12440 19728 12492 19780
rect 12992 19728 13044 19780
rect 20444 19771 20496 19780
rect 20444 19737 20453 19771
rect 20453 19737 20487 19771
rect 20487 19737 20496 19771
rect 20444 19728 20496 19737
rect 57060 19864 57112 19916
rect 57796 19907 57848 19916
rect 57796 19873 57805 19907
rect 57805 19873 57839 19907
rect 57839 19873 57848 19907
rect 57796 19864 57848 19873
rect 46756 19728 46808 19780
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 2504 19499 2556 19508
rect 2504 19465 2513 19499
rect 2513 19465 2547 19499
rect 2547 19465 2556 19499
rect 2504 19456 2556 19465
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 12440 19320 12492 19372
rect 19432 19320 19484 19372
rect 20076 19363 20128 19372
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20076 19320 20128 19329
rect 29644 19320 29696 19372
rect 30380 19320 30432 19372
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2228 18708 2280 18760
rect 9036 18708 9088 18760
rect 2412 18572 2464 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2412 18343 2464 18352
rect 2412 18309 2421 18343
rect 2421 18309 2455 18343
rect 2455 18309 2464 18343
rect 2412 18300 2464 18309
rect 2228 18275 2280 18284
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 30380 18275 30432 18284
rect 30380 18241 30389 18275
rect 30389 18241 30423 18275
rect 30423 18241 30432 18275
rect 30380 18232 30432 18241
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 31208 18028 31260 18080
rect 56876 18028 56928 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 31024 17731 31076 17740
rect 31024 17697 31033 17731
rect 31033 17697 31067 17731
rect 31067 17697 31076 17731
rect 31024 17688 31076 17697
rect 31208 17731 31260 17740
rect 31208 17697 31217 17731
rect 31217 17697 31251 17731
rect 31251 17697 31260 17731
rect 31208 17688 31260 17697
rect 56876 17688 56928 17740
rect 58164 17731 58216 17740
rect 58164 17697 58173 17731
rect 58173 17697 58207 17731
rect 58207 17697 58216 17731
rect 58164 17688 58216 17697
rect 1952 17620 2004 17672
rect 32864 17595 32916 17604
rect 32864 17561 32873 17595
rect 32873 17561 32907 17595
rect 32907 17561 32916 17595
rect 32864 17552 32916 17561
rect 57152 17552 57204 17604
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 57152 17323 57204 17332
rect 57152 17289 57161 17323
rect 57161 17289 57195 17323
rect 57195 17289 57204 17323
rect 57152 17280 57204 17289
rect 1952 17187 2004 17196
rect 1952 17153 1961 17187
rect 1961 17153 1995 17187
rect 1995 17153 2004 17187
rect 1952 17144 2004 17153
rect 17408 17144 17460 17196
rect 20076 17144 20128 17196
rect 57060 17187 57112 17196
rect 57060 17153 57069 17187
rect 57069 17153 57103 17187
rect 57103 17153 57112 17187
rect 57060 17144 57112 17153
rect 2136 17119 2188 17128
rect 2136 17085 2145 17119
rect 2145 17085 2179 17119
rect 2179 17085 2188 17119
rect 2136 17076 2188 17085
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 56324 16940 56376 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2136 16736 2188 16788
rect 2044 16600 2096 16652
rect 29552 16600 29604 16652
rect 30288 16600 30340 16652
rect 56324 16643 56376 16652
rect 56324 16609 56333 16643
rect 56333 16609 56367 16643
rect 56367 16609 56376 16643
rect 56324 16600 56376 16609
rect 57796 16643 57848 16652
rect 57796 16609 57805 16643
rect 57805 16609 57839 16643
rect 57839 16609 57848 16643
rect 57796 16600 57848 16609
rect 57152 16464 57204 16516
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 57152 16235 57204 16244
rect 57152 16201 57161 16235
rect 57161 16201 57195 16235
rect 57195 16201 57204 16235
rect 57152 16192 57204 16201
rect 57060 16099 57112 16108
rect 57060 16065 57069 16099
rect 57069 16065 57103 16099
rect 57103 16065 57112 16099
rect 57060 16056 57112 16065
rect 56324 15852 56376 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 56324 15555 56376 15564
rect 56324 15521 56333 15555
rect 56333 15521 56367 15555
rect 56367 15521 56376 15555
rect 56324 15512 56376 15521
rect 57888 15555 57940 15564
rect 57888 15521 57897 15555
rect 57897 15521 57931 15555
rect 57931 15521 57940 15555
rect 57888 15512 57940 15521
rect 56968 15376 57020 15428
rect 57060 15308 57112 15360
rect 57796 15308 57848 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 56968 15147 57020 15156
rect 56968 15113 56977 15147
rect 56977 15113 57011 15147
rect 57011 15113 57020 15147
rect 56968 15104 57020 15113
rect 55680 14968 55732 15020
rect 57336 14968 57388 15020
rect 56324 14764 56376 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 56324 14467 56376 14476
rect 56324 14433 56333 14467
rect 56333 14433 56367 14467
rect 56367 14433 56376 14467
rect 56324 14424 56376 14433
rect 1952 14356 2004 14408
rect 56968 14288 57020 14340
rect 58164 14331 58216 14340
rect 58164 14297 58173 14331
rect 58173 14297 58207 14331
rect 58207 14297 58216 14331
rect 58164 14288 58216 14297
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 56968 14059 57020 14068
rect 56968 14025 56977 14059
rect 56977 14025 57011 14059
rect 57011 14025 57020 14059
rect 56968 14016 57020 14025
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 57152 13880 57204 13932
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2136 13472 2188 13524
rect 2688 13268 2740 13320
rect 4712 13268 4764 13320
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 3884 12724 3936 12776
rect 3976 12767 4028 12776
rect 3976 12733 3985 12767
rect 3985 12733 4019 12767
rect 4019 12733 4028 12767
rect 3976 12724 4028 12733
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 1952 12180 2004 12232
rect 14832 12180 14884 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2412 11636 2464 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2412 11339 2464 11348
rect 2412 11305 2421 11339
rect 2421 11305 2455 11339
rect 2455 11305 2464 11339
rect 2412 11296 2464 11305
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 9128 11092 9180 11144
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 20352 10140 20404 10192
rect 56692 10140 56744 10192
rect 3424 9936 3476 9988
rect 29368 10004 29420 10056
rect 29736 9979 29788 9988
rect 29736 9945 29745 9979
rect 29745 9945 29779 9979
rect 29779 9945 29788 9979
rect 29736 9936 29788 9945
rect 27160 9868 27212 9920
rect 56692 10004 56744 10056
rect 57244 9979 57296 9988
rect 57244 9945 57253 9979
rect 57253 9945 57287 9979
rect 57287 9945 57296 9979
rect 57244 9936 57296 9945
rect 56692 9911 56744 9920
rect 56692 9877 56701 9911
rect 56701 9877 56735 9911
rect 56735 9877 56744 9911
rect 56692 9868 56744 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 29736 9664 29788 9716
rect 29552 9571 29604 9580
rect 29552 9537 29561 9571
rect 29561 9537 29595 9571
rect 29595 9537 29604 9571
rect 29552 9528 29604 9537
rect 56324 9324 56376 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 56324 9027 56376 9036
rect 56324 8993 56333 9027
rect 56333 8993 56367 9027
rect 56367 8993 56376 9027
rect 56324 8984 56376 8993
rect 56692 8984 56744 9036
rect 57888 9027 57940 9036
rect 57888 8993 57897 9027
rect 57897 8993 57931 9027
rect 57931 8993 57940 9027
rect 57888 8984 57940 8993
rect 1952 8916 2004 8968
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 1952 7828 2004 7880
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 9864 7828 9916 7880
rect 2136 7692 2188 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 2136 7463 2188 7472
rect 2136 7429 2145 7463
rect 2145 7429 2179 7463
rect 2179 7429 2188 7463
rect 2136 7420 2188 7429
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 20260 7352 20312 7404
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 4620 7148 4672 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4620 6740 4672 6792
rect 20444 6740 20496 6792
rect 56876 6740 56928 6792
rect 3240 6715 3292 6724
rect 3240 6681 3249 6715
rect 3249 6681 3283 6715
rect 3283 6681 3292 6715
rect 3240 6672 3292 6681
rect 56324 6672 56376 6724
rect 57060 6647 57112 6656
rect 57060 6613 57069 6647
rect 57069 6613 57103 6647
rect 57103 6613 57112 6647
rect 57060 6604 57112 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 2964 6332 3016 6384
rect 5172 6375 5224 6384
rect 5172 6341 5181 6375
rect 5181 6341 5215 6375
rect 5215 6341 5224 6375
rect 5172 6332 5224 6341
rect 7840 6332 7892 6384
rect 29460 6264 29512 6316
rect 1860 6196 1912 6248
rect 2412 6196 2464 6248
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 56600 6060 56652 6112
rect 57336 6060 57388 6112
rect 57980 6103 58032 6112
rect 57980 6069 57989 6103
rect 57989 6069 58023 6103
rect 58023 6069 58032 6103
rect 57980 6060 58032 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 56324 5763 56376 5772
rect 56324 5729 56333 5763
rect 56333 5729 56367 5763
rect 56367 5729 56376 5763
rect 56324 5720 56376 5729
rect 57980 5720 58032 5772
rect 58164 5763 58216 5772
rect 58164 5729 58173 5763
rect 58173 5729 58207 5763
rect 58207 5729 58216 5763
rect 58164 5720 58216 5729
rect 2044 5652 2096 5704
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 55496 5652 55548 5704
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 3056 5244 3108 5296
rect 57060 5244 57112 5296
rect 55496 5219 55548 5228
rect 55496 5185 55505 5219
rect 55505 5185 55539 5219
rect 55539 5185 55548 5219
rect 55496 5176 55548 5185
rect 1860 5108 1912 5160
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 58624 5108 58676 5160
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 56324 4972 56376 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 56324 4675 56376 4684
rect 56324 4641 56333 4675
rect 56333 4641 56367 4675
rect 56367 4641 56376 4675
rect 56324 4632 56376 4641
rect 56508 4632 56560 4684
rect 2228 4564 2280 4616
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 22836 4564 22888 4616
rect 55036 4564 55088 4616
rect 55496 4564 55548 4616
rect 57980 4496 58032 4548
rect 8208 4428 8260 4480
rect 9588 4428 9640 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 8208 4199 8260 4208
rect 8208 4165 8217 4199
rect 8217 4165 8251 4199
rect 8251 4165 8260 4199
rect 8208 4156 8260 4165
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 14832 4131 14884 4140
rect 1860 4020 1912 4072
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 2780 4020 2832 4029
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 22468 4131 22520 4140
rect 14832 4088 14884 4097
rect 8300 4020 8352 4072
rect 8392 4020 8444 4072
rect 22468 4097 22477 4131
rect 22477 4097 22511 4131
rect 22511 4097 22520 4131
rect 22468 4088 22520 4097
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 29828 4088 29880 4140
rect 31116 4131 31168 4140
rect 31116 4097 31125 4131
rect 31125 4097 31159 4131
rect 31159 4097 31168 4131
rect 31116 4088 31168 4097
rect 49976 4131 50028 4140
rect 29184 4020 29236 4072
rect 30564 3952 30616 4004
rect 49976 4097 49985 4131
rect 49985 4097 50019 4131
rect 50019 4097 50028 4131
rect 49976 4088 50028 4097
rect 53840 4131 53892 4140
rect 53840 4097 53849 4131
rect 53849 4097 53883 4131
rect 53883 4097 53892 4131
rect 53840 4088 53892 4097
rect 56600 4156 56652 4208
rect 55496 4131 55548 4140
rect 46756 4020 46808 4072
rect 55496 4097 55505 4131
rect 55505 4097 55539 4131
rect 55539 4097 55548 4131
rect 55496 4088 55548 4097
rect 57796 4088 57848 4140
rect 44548 3952 44600 4004
rect 57704 4020 57756 4072
rect 3792 3884 3844 3936
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 15292 3884 15344 3936
rect 16672 3884 16724 3936
rect 23020 3884 23072 3936
rect 23296 3927 23348 3936
rect 23296 3893 23305 3927
rect 23305 3893 23339 3927
rect 23339 3893 23348 3927
rect 23296 3884 23348 3893
rect 26884 3884 26936 3936
rect 29736 3884 29788 3936
rect 30656 3927 30708 3936
rect 30656 3893 30665 3927
rect 30665 3893 30699 3927
rect 30699 3893 30708 3927
rect 30656 3884 30708 3893
rect 30748 3884 30800 3936
rect 32128 3884 32180 3936
rect 38476 3884 38528 3936
rect 46296 3884 46348 3936
rect 50344 3884 50396 3936
rect 53104 3884 53156 3936
rect 55404 3884 55456 3936
rect 57152 3884 57204 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 1860 3723 1912 3732
rect 1860 3689 1869 3723
rect 1869 3689 1903 3723
rect 1903 3689 1912 3723
rect 1860 3680 1912 3689
rect 8944 3680 8996 3732
rect 22468 3680 22520 3732
rect 56784 3680 56836 3732
rect 3792 3587 3844 3596
rect 3792 3553 3801 3587
rect 3801 3553 3835 3587
rect 3835 3553 3844 3587
rect 3792 3544 3844 3553
rect 3976 3544 4028 3596
rect 5172 3544 5224 3596
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 9680 3544 9732 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 2320 3340 2372 3392
rect 5356 3476 5408 3528
rect 12256 3519 12308 3528
rect 6276 3451 6328 3460
rect 6276 3417 6285 3451
rect 6285 3417 6319 3451
rect 6319 3417 6328 3451
rect 6276 3408 6328 3417
rect 12256 3485 12265 3519
rect 12265 3485 12299 3519
rect 12299 3485 12308 3519
rect 12256 3476 12308 3485
rect 12532 3476 12584 3528
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 9772 3408 9824 3460
rect 15476 3408 15528 3460
rect 9220 3340 9272 3392
rect 12716 3340 12768 3392
rect 16856 3340 16908 3392
rect 32956 3612 33008 3664
rect 43260 3612 43312 3664
rect 20628 3544 20680 3596
rect 25136 3587 25188 3596
rect 25136 3553 25145 3587
rect 25145 3553 25179 3587
rect 25179 3553 25188 3587
rect 25136 3544 25188 3553
rect 26884 3587 26936 3596
rect 26884 3553 26893 3587
rect 26893 3553 26927 3587
rect 26927 3553 26936 3587
rect 26884 3544 26936 3553
rect 27068 3544 27120 3596
rect 30656 3544 30708 3596
rect 32128 3587 32180 3596
rect 32128 3553 32137 3587
rect 32137 3553 32171 3587
rect 32171 3553 32180 3587
rect 32128 3544 32180 3553
rect 32864 3587 32916 3596
rect 32864 3553 32873 3587
rect 32873 3553 32907 3587
rect 32907 3553 32916 3587
rect 32864 3544 32916 3553
rect 34152 3544 34204 3596
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 22836 3519 22888 3528
rect 22836 3485 22845 3519
rect 22845 3485 22879 3519
rect 22879 3485 22888 3519
rect 22836 3476 22888 3485
rect 26700 3519 26752 3528
rect 26700 3485 26709 3519
rect 26709 3485 26743 3519
rect 26743 3485 26752 3519
rect 26700 3476 26752 3485
rect 38292 3476 38344 3528
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 47032 3587 47084 3596
rect 47032 3553 47041 3587
rect 47041 3553 47075 3587
rect 47075 3553 47084 3587
rect 47032 3544 47084 3553
rect 50344 3587 50396 3596
rect 50344 3553 50353 3587
rect 50353 3553 50387 3587
rect 50387 3553 50396 3587
rect 50344 3544 50396 3553
rect 50620 3587 50672 3596
rect 50620 3553 50629 3587
rect 50629 3553 50663 3587
rect 50663 3553 50672 3587
rect 50620 3544 50672 3553
rect 53104 3587 53156 3596
rect 53104 3553 53113 3587
rect 53113 3553 53147 3587
rect 53147 3553 53156 3587
rect 53104 3544 53156 3553
rect 54116 3587 54168 3596
rect 54116 3553 54125 3587
rect 54125 3553 54159 3587
rect 54159 3553 54168 3587
rect 54116 3544 54168 3553
rect 48228 3476 48280 3528
rect 52920 3519 52972 3528
rect 52920 3485 52929 3519
rect 52929 3485 52963 3519
rect 52963 3485 52972 3519
rect 52920 3476 52972 3485
rect 28816 3408 28868 3460
rect 31208 3408 31260 3460
rect 31576 3408 31628 3460
rect 32680 3408 32732 3460
rect 43260 3408 43312 3460
rect 26976 3340 27028 3392
rect 44548 3340 44600 3392
rect 46848 3408 46900 3460
rect 57612 3612 57664 3664
rect 57888 3587 57940 3596
rect 57888 3553 57897 3587
rect 57897 3553 57931 3587
rect 57931 3553 57940 3587
rect 57888 3544 57940 3553
rect 58072 3476 58124 3528
rect 56048 3408 56100 3460
rect 56968 3408 57020 3460
rect 48320 3340 48372 3392
rect 54208 3340 54260 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 6276 3136 6328 3188
rect 2320 3111 2372 3120
rect 2320 3077 2329 3111
rect 2329 3077 2363 3111
rect 2363 3077 2372 3111
rect 2320 3068 2372 3077
rect 12256 3068 12308 3120
rect 12716 3111 12768 3120
rect 12716 3077 12725 3111
rect 12725 3077 12759 3111
rect 12759 3077 12768 3111
rect 12716 3068 12768 3077
rect 16856 3111 16908 3120
rect 16856 3077 16865 3111
rect 16865 3077 16899 3111
rect 16899 3077 16908 3111
rect 16856 3068 16908 3077
rect 4712 3000 4764 3052
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 15108 3000 15160 3052
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 20352 3000 20404 3052
rect 23296 3136 23348 3188
rect 32680 3179 32732 3188
rect 32680 3145 32689 3179
rect 32689 3145 32723 3179
rect 32723 3145 32732 3179
rect 32680 3136 32732 3145
rect 46848 3179 46900 3188
rect 46848 3145 46857 3179
rect 46857 3145 46891 3179
rect 46891 3145 46900 3179
rect 46848 3136 46900 3145
rect 49976 3136 50028 3188
rect 56968 3179 57020 3188
rect 23020 3111 23072 3120
rect 23020 3077 23029 3111
rect 23029 3077 23063 3111
rect 23063 3077 23072 3111
rect 23020 3068 23072 3077
rect 30748 3068 30800 3120
rect 38476 3111 38528 3120
rect 38476 3077 38485 3111
rect 38485 3077 38519 3111
rect 38519 3077 38528 3111
rect 38476 3068 38528 3077
rect 54208 3111 54260 3120
rect 54208 3077 54217 3111
rect 54217 3077 54251 3111
rect 54251 3077 54260 3111
rect 54208 3068 54260 3077
rect 56968 3145 56977 3179
rect 56977 3145 57011 3179
rect 57011 3145 57020 3179
rect 56968 3136 57020 3145
rect 57980 3179 58032 3188
rect 57980 3145 57989 3179
rect 57989 3145 58023 3179
rect 58023 3145 58032 3179
rect 57980 3136 58032 3145
rect 26700 3000 26752 3052
rect 29736 3043 29788 3052
rect 29736 3009 29745 3043
rect 29745 3009 29779 3043
rect 29779 3009 29788 3043
rect 29736 3000 29788 3009
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 664 2864 716 2916
rect 9036 2932 9088 2984
rect 7748 2864 7800 2916
rect 12900 2932 12952 2984
rect 16120 2932 16172 2984
rect 23204 2932 23256 2984
rect 30932 2975 30984 2984
rect 30932 2941 30941 2975
rect 30941 2941 30975 2975
rect 30975 2941 30984 2975
rect 30932 2932 30984 2941
rect 38292 3043 38344 3052
rect 38292 3009 38301 3043
rect 38301 3009 38335 3043
rect 38335 3009 38344 3043
rect 38292 3000 38344 3009
rect 46756 3043 46808 3052
rect 46756 3009 46765 3043
rect 46765 3009 46799 3043
rect 46799 3009 46808 3043
rect 46756 3000 46808 3009
rect 47584 3043 47636 3052
rect 47584 3009 47593 3043
rect 47593 3009 47627 3043
rect 47627 3009 47636 3043
rect 47584 3000 47636 3009
rect 48228 3043 48280 3052
rect 48228 3009 48237 3043
rect 48237 3009 48271 3043
rect 48271 3009 48280 3043
rect 48228 3000 48280 3009
rect 52920 3000 52972 3052
rect 56784 3000 56836 3052
rect 38660 2932 38712 2984
rect 49608 2975 49660 2984
rect 49608 2941 49617 2975
rect 49617 2941 49651 2975
rect 49651 2941 49660 2975
rect 49608 2932 49660 2941
rect 54024 2975 54076 2984
rect 54024 2941 54033 2975
rect 54033 2941 54067 2975
rect 54067 2941 54076 2975
rect 54024 2932 54076 2941
rect 54760 2975 54812 2984
rect 54760 2941 54769 2975
rect 54769 2941 54803 2975
rect 54803 2941 54812 2975
rect 54760 2932 54812 2941
rect 6920 2839 6972 2848
rect 6920 2805 6929 2839
rect 6929 2805 6963 2839
rect 6963 2805 6972 2839
rect 6920 2796 6972 2805
rect 28816 2796 28868 2848
rect 31116 2796 31168 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2136 2592 2188 2644
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 31208 2635 31260 2644
rect 31208 2601 31217 2635
rect 31217 2601 31251 2635
rect 31251 2601 31260 2635
rect 31208 2592 31260 2601
rect 54024 2592 54076 2644
rect 58072 2635 58124 2644
rect 58072 2601 58081 2635
rect 58081 2601 58115 2635
rect 58115 2601 58124 2635
rect 58072 2592 58124 2601
rect 6460 2524 6512 2576
rect 6920 2456 6972 2508
rect 53840 2456 53892 2508
rect 55036 2456 55088 2508
rect 31116 2431 31168 2440
rect 31116 2397 31125 2431
rect 31125 2397 31159 2431
rect 31159 2397 31168 2431
rect 31116 2388 31168 2397
rect 7472 2320 7524 2372
rect 55404 2320 55456 2372
rect 57336 2363 57388 2372
rect 57336 2329 57345 2363
rect 57345 2329 57379 2363
rect 57379 2329 57388 2363
rect 57336 2320 57388 2329
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 634 59200 746 60000
rect 1278 59200 1390 60000
rect 2566 59200 2678 60000
rect 3854 59200 3966 60000
rect 5142 59200 5254 60000
rect 5786 59200 5898 60000
rect 7074 59200 7186 60000
rect 8362 59200 8474 60000
rect 9650 59200 9762 60000
rect 10294 59200 10406 60000
rect 11582 59200 11694 60000
rect 12870 59200 12982 60000
rect 13514 59200 13626 60000
rect 14802 59200 14914 60000
rect 16090 59200 16202 60000
rect 17378 59200 17490 60000
rect 18022 59200 18134 60000
rect 19310 59200 19422 60000
rect 20598 59200 20710 60000
rect 21242 59200 21354 60000
rect 22530 59200 22642 60000
rect 23818 59200 23930 60000
rect 25106 59200 25218 60000
rect 25750 59200 25862 60000
rect 27038 59200 27150 60000
rect 28326 59200 28438 60000
rect 28970 59200 29082 60000
rect 30258 59200 30370 60000
rect 31546 59200 31658 60000
rect 32834 59200 32946 60000
rect 33478 59200 33590 60000
rect 34766 59200 34878 60000
rect 36054 59200 36166 60000
rect 36698 59200 36810 60000
rect 37986 59200 38098 60000
rect 39274 59200 39386 60000
rect 40562 59200 40674 60000
rect 41206 59200 41318 60000
rect 42494 59200 42606 60000
rect 43782 59200 43894 60000
rect 44426 59200 44538 60000
rect 45714 59200 45826 60000
rect 47002 59200 47114 60000
rect 48290 59200 48402 60000
rect 48934 59200 49046 60000
rect 50222 59200 50334 60000
rect 51510 59200 51622 60000
rect 52154 59200 52266 60000
rect 53442 59200 53554 60000
rect 54730 59200 54842 60000
rect 56018 59200 56130 60000
rect 56662 59200 56774 60000
rect 57950 59200 58062 60000
rect 59238 59200 59350 60000
rect 59882 59200 59994 60000
rect 676 57458 704 59200
rect 664 57452 716 57458
rect 664 57394 716 57400
rect 1952 56840 2004 56846
rect 1952 56782 2004 56788
rect 1964 56370 1992 56782
rect 1952 56364 2004 56370
rect 1952 56306 2004 56312
rect 2136 56296 2188 56302
rect 2136 56238 2188 56244
rect 1490 55856 1546 55865
rect 1490 55791 1546 55800
rect 1504 55758 1532 55791
rect 1492 55752 1544 55758
rect 1492 55694 1544 55700
rect 2044 55684 2096 55690
rect 2044 55626 2096 55632
rect 1952 53576 2004 53582
rect 1952 53518 2004 53524
rect 1964 53106 1992 53518
rect 1952 53100 2004 53106
rect 1952 53042 2004 53048
rect 2056 45558 2084 55626
rect 2148 54874 2176 56238
rect 2608 55622 2636 59200
rect 2778 57896 2834 57905
rect 2778 57831 2834 57840
rect 2792 56302 2820 57831
rect 3896 57610 3924 59200
rect 3896 57582 4108 57610
rect 3700 57248 3752 57254
rect 3700 57190 3752 57196
rect 3792 57248 3844 57254
rect 3792 57190 3844 57196
rect 3974 57216 4030 57225
rect 2872 56840 2924 56846
rect 2872 56782 2924 56788
rect 2780 56296 2832 56302
rect 2780 56238 2832 56244
rect 2596 55616 2648 55622
rect 2596 55558 2648 55564
rect 2884 55350 2912 56782
rect 3712 55758 3740 57190
rect 3804 56914 3832 57190
rect 3974 57151 4030 57160
rect 3792 56908 3844 56914
rect 3792 56850 3844 56856
rect 3700 55752 3752 55758
rect 3700 55694 3752 55700
rect 2872 55344 2924 55350
rect 2872 55286 2924 55292
rect 3988 55214 4016 57151
rect 4080 56930 4108 57582
rect 4214 57148 4522 57168
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57072 4522 57092
rect 4080 56914 4200 56930
rect 4080 56908 4212 56914
rect 4080 56902 4160 56908
rect 4160 56850 4212 56856
rect 4344 56772 4396 56778
rect 4344 56714 4396 56720
rect 4356 56506 4384 56714
rect 4344 56500 4396 56506
rect 4344 56442 4396 56448
rect 5828 56234 5856 59200
rect 6368 56840 6420 56846
rect 6368 56782 6420 56788
rect 6380 56370 6408 56782
rect 6368 56364 6420 56370
rect 6368 56306 6420 56312
rect 6920 56296 6972 56302
rect 6920 56238 6972 56244
rect 5816 56228 5868 56234
rect 5816 56170 5868 56176
rect 4712 56160 4764 56166
rect 4712 56102 4764 56108
rect 4214 56060 4522 56080
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55984 4522 56004
rect 3792 55208 3844 55214
rect 3792 55150 3844 55156
rect 3976 55208 4028 55214
rect 3976 55150 4028 55156
rect 3804 54874 3832 55150
rect 4214 54972 4522 54992
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54896 4522 54916
rect 2136 54868 2188 54874
rect 2136 54810 2188 54816
rect 3792 54868 3844 54874
rect 3792 54810 3844 54816
rect 3332 54664 3384 54670
rect 3332 54606 3384 54612
rect 3976 54664 4028 54670
rect 3976 54606 4028 54612
rect 2778 54496 2834 54505
rect 2778 54431 2834 54440
rect 2792 53038 2820 54431
rect 2412 53032 2464 53038
rect 2412 52974 2464 52980
rect 2780 53032 2832 53038
rect 2780 52974 2832 52980
rect 2424 52698 2452 52974
rect 2412 52692 2464 52698
rect 2412 52634 2464 52640
rect 2320 52488 2372 52494
rect 2320 52430 2372 52436
rect 3148 52488 3200 52494
rect 3148 52430 3200 52436
rect 3238 52456 3294 52465
rect 2044 45552 2096 45558
rect 2044 45494 2096 45500
rect 2056 44470 2084 45494
rect 2044 44464 2096 44470
rect 2044 44406 2096 44412
rect 2228 39840 2280 39846
rect 2228 39782 2280 39788
rect 2240 38962 2268 39782
rect 2228 38956 2280 38962
rect 2228 38898 2280 38904
rect 1952 30048 2004 30054
rect 1952 29990 2004 29996
rect 2136 30048 2188 30054
rect 2136 29990 2188 29996
rect 1964 29170 1992 29990
rect 2148 29238 2176 29990
rect 2136 29232 2188 29238
rect 2136 29174 2188 29180
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 1964 26994 1992 27406
rect 1952 26988 2004 26994
rect 1952 26930 2004 26936
rect 2332 24818 2360 52430
rect 3160 51950 3188 52430
rect 3238 52391 3294 52400
rect 3252 51950 3280 52391
rect 3148 51944 3200 51950
rect 3148 51886 3200 51892
rect 3240 51944 3292 51950
rect 3240 51886 3292 51892
rect 2962 49056 3018 49065
rect 2962 48991 3018 49000
rect 2976 47258 3004 48991
rect 2964 47252 3016 47258
rect 2964 47194 3016 47200
rect 3344 45554 3372 54606
rect 3884 52352 3936 52358
rect 3884 52294 3936 52300
rect 3896 52086 3924 52294
rect 3884 52080 3936 52086
rect 3884 52022 3936 52028
rect 3424 49768 3476 49774
rect 3422 49736 3424 49745
rect 3476 49736 3478 49745
rect 3422 49671 3478 49680
rect 3344 45526 3464 45554
rect 3436 45014 3464 45526
rect 3424 45008 3476 45014
rect 3424 44950 3476 44956
rect 2688 44464 2740 44470
rect 2688 44406 2740 44412
rect 2412 39296 2464 39302
rect 2412 39238 2464 39244
rect 2424 39030 2452 39238
rect 2412 39024 2464 39030
rect 2412 38966 2464 38972
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 1964 23730 1992 24550
rect 2148 23798 2176 24550
rect 2136 23792 2188 23798
rect 2136 23734 2188 23740
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1964 21554 1992 21966
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1964 20466 1992 20878
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 2148 20058 2176 21422
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2240 18290 2268 18702
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1964 17202 1992 17614
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2148 16794 2176 17070
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 13938 1992 14350
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1964 11762 1992 12174
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1964 8498 1992 8910
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2056 7886 2084 16594
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2148 13530 2176 13806
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2332 11150 2360 24754
rect 2424 19378 2452 30194
rect 2504 26920 2556 26926
rect 2504 26862 2556 26868
rect 2516 26586 2544 26862
rect 2504 26580 2556 26586
rect 2504 26522 2556 26528
rect 2700 25974 2728 44406
rect 3436 44198 3464 44950
rect 2964 44192 3016 44198
rect 2964 44134 3016 44140
rect 3424 44192 3476 44198
rect 3424 44134 3476 44140
rect 2778 39536 2834 39545
rect 2778 39471 2834 39480
rect 2792 38894 2820 39471
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 2778 30016 2834 30025
rect 2778 29951 2834 29960
rect 2792 29102 2820 29951
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2792 26625 2820 26862
rect 2778 26616 2834 26625
rect 2778 26551 2834 26560
rect 2688 25968 2740 25974
rect 2688 25910 2740 25916
rect 2778 24576 2834 24585
rect 2778 24511 2834 24520
rect 2792 23662 2820 24511
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2778 21856 2834 21865
rect 2778 21791 2834 21800
rect 2792 21486 2820 21791
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2778 20496 2834 20505
rect 2778 20431 2834 20440
rect 2792 20398 2820 20431
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2516 19514 2544 20334
rect 2688 19848 2740 19854
rect 2688 19790 2740 19796
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2412 18624 2464 18630
rect 2412 18566 2464 18572
rect 2424 18358 2452 18566
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2700 13326 2728 19790
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 18222 2820 18391
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2780 17128 2832 17134
rect 2778 17096 2780 17105
rect 2832 17096 2834 17105
rect 2778 17031 2834 17040
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13705 2820 13806
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2412 11688 2464 11694
rect 2780 11688 2832 11694
rect 2412 11630 2464 11636
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2424 11354 2452 11630
rect 2778 11591 2834 11600
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2148 8090 2176 8366
rect 2792 8265 2820 8366
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 1964 7410 1992 7822
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 5914 1900 6190
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2056 5710 2084 7822
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2148 7478 2176 7686
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2792 6905 2820 7278
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2976 6390 3004 44134
rect 3884 39432 3936 39438
rect 3884 39374 3936 39380
rect 3424 29028 3476 29034
rect 3424 28970 3476 28976
rect 3436 28665 3464 28970
rect 3422 28656 3478 28665
rect 3422 28591 3478 28600
rect 3896 21350 3924 39374
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3988 20398 4016 54606
rect 4214 53884 4522 53904
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53808 4522 53828
rect 4214 52796 4522 52816
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52720 4522 52740
rect 4214 51708 4522 51728
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51632 4522 51652
rect 4214 50620 4522 50640
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50544 4522 50564
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4724 45554 4752 56102
rect 6932 55962 6960 56238
rect 7116 56234 7144 59200
rect 10336 57458 10364 59200
rect 10324 57452 10376 57458
rect 10324 57394 10376 57400
rect 8668 56840 8720 56846
rect 8668 56782 8720 56788
rect 13268 56840 13320 56846
rect 13268 56782 13320 56788
rect 8680 56370 8708 56782
rect 13280 56370 13308 56782
rect 8668 56364 8720 56370
rect 8668 56306 8720 56312
rect 13268 56364 13320 56370
rect 13268 56306 13320 56312
rect 13556 56302 13584 59200
rect 16028 56840 16080 56846
rect 16028 56782 16080 56788
rect 9036 56296 9088 56302
rect 9036 56238 9088 56244
rect 13084 56296 13136 56302
rect 13084 56238 13136 56244
rect 13544 56296 13596 56302
rect 13544 56238 13596 56244
rect 7104 56228 7156 56234
rect 7104 56170 7156 56176
rect 9048 55962 9076 56238
rect 13096 55962 13124 56238
rect 15108 56160 15160 56166
rect 15108 56102 15160 56108
rect 6920 55956 6972 55962
rect 6920 55898 6972 55904
rect 9036 55956 9088 55962
rect 9036 55898 9088 55904
rect 13084 55956 13136 55962
rect 13084 55898 13136 55904
rect 9496 55888 9548 55894
rect 9496 55830 9548 55836
rect 8944 55752 8996 55758
rect 8944 55694 8996 55700
rect 5172 53168 5224 53174
rect 5172 53110 5224 53116
rect 5184 52494 5212 53110
rect 5172 52488 5224 52494
rect 5172 52430 5224 52436
rect 4632 45526 4752 45554
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4632 39438 4660 45526
rect 4620 39432 4672 39438
rect 4620 39374 4672 39380
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3896 12442 3924 12718
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3988 12345 4016 12718
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3974 12336 4030 12345
rect 3974 12271 4030 12280
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3436 8945 3464 9930
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 3422 8936 3478 8945
rect 3422 8871 3478 8880
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4632 6798 4660 7142
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2424 5914 2452 6190
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 1872 4826 1900 5102
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2240 4146 2268 4558
rect 2792 4185 2820 5102
rect 2778 4176 2834 4185
rect 2228 4140 2280 4146
rect 2778 4111 2834 4120
rect 2228 4082 2280 4088
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 1872 3738 1900 4014
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3126 2360 3334
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 676 800 704 2858
rect 2148 2650 2176 2926
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2792 2145 2820 4014
rect 2884 3505 2912 6190
rect 2976 5710 3004 6326
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3056 5568 3108 5574
rect 3252 5545 3280 6666
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3056 5510 3108 5516
rect 3238 5536 3294 5545
rect 3068 5302 3096 5510
rect 3238 5471 3294 5480
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3602 3832 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 3988 1714 4016 3538
rect 4724 3058 4752 13262
rect 5184 6390 5212 52430
rect 8484 48680 8536 48686
rect 8484 48622 8536 48628
rect 8496 27130 8524 48622
rect 8956 47666 8984 55694
rect 8944 47660 8996 47666
rect 8944 47602 8996 47608
rect 8484 27124 8536 27130
rect 8484 27066 8536 27072
rect 8760 26988 8812 26994
rect 8760 26930 8812 26936
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8588 24818 8616 26862
rect 8772 26382 8800 26930
rect 8760 26376 8812 26382
rect 8760 26318 8812 26324
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 8772 25906 8800 26318
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8772 25294 8800 25842
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8772 24818 8800 25230
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 9036 24744 9088 24750
rect 9036 24686 9088 24692
rect 9048 18766 9076 24686
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 9048 6914 9076 18702
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8956 6886 9076 6914
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7852 4622 7880 6326
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4214 8248 4422
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8312 4078 8340 4966
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3896 1686 4016 1714
rect 3896 800 3924 1686
rect 5184 800 5212 3538
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5368 3058 5396 3470
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 6288 3194 6316 3402
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 6472 800 6500 2518
rect 6932 2514 6960 2790
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7484 2378 7512 3878
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7760 800 7788 2858
rect 8404 800 8432 4014
rect 8956 3738 8984 6886
rect 9140 4622 9168 11086
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9232 3398 9260 26318
rect 9508 25838 9536 55830
rect 15120 55758 15148 56102
rect 16040 55826 16068 56782
rect 16132 55826 16160 59200
rect 17316 56840 17368 56846
rect 17316 56782 17368 56788
rect 17132 56296 17184 56302
rect 17132 56238 17184 56244
rect 16028 55820 16080 55826
rect 16028 55762 16080 55768
rect 16120 55820 16172 55826
rect 16120 55762 16172 55768
rect 12992 55752 13044 55758
rect 12992 55694 13044 55700
rect 15108 55752 15160 55758
rect 15108 55694 15160 55700
rect 9680 49768 9732 49774
rect 9680 49710 9732 49716
rect 9692 48686 9720 49710
rect 9680 48680 9732 48686
rect 9680 48622 9732 48628
rect 9864 25968 9916 25974
rect 9864 25910 9916 25916
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9876 25226 9904 25910
rect 9864 25220 9916 25226
rect 9864 25162 9916 25168
rect 9876 7886 9904 25162
rect 13004 19786 13032 55694
rect 16580 55616 16632 55622
rect 16580 55558 16632 55564
rect 16592 25974 16620 55558
rect 16580 25968 16632 25974
rect 16580 25910 16632 25916
rect 17144 21690 17172 56238
rect 17328 55622 17356 56782
rect 17420 56302 17448 59200
rect 18064 57254 18092 59200
rect 17960 57248 18012 57254
rect 17960 57190 18012 57196
rect 18052 57248 18104 57254
rect 18052 57190 18104 57196
rect 19248 57248 19300 57254
rect 19248 57190 19300 57196
rect 17868 56704 17920 56710
rect 17868 56646 17920 56652
rect 17408 56296 17460 56302
rect 17408 56238 17460 56244
rect 17316 55616 17368 55622
rect 17316 55558 17368 55564
rect 17880 55214 17908 56646
rect 17972 55350 18000 57190
rect 18236 56840 18288 56846
rect 18236 56782 18288 56788
rect 18248 56438 18276 56782
rect 18236 56432 18288 56438
rect 18236 56374 18288 56380
rect 19064 56296 19116 56302
rect 19064 56238 19116 56244
rect 19076 55894 19104 56238
rect 19064 55888 19116 55894
rect 19064 55830 19116 55836
rect 17960 55344 18012 55350
rect 17960 55286 18012 55292
rect 19260 55214 19288 57190
rect 19352 56302 19380 59200
rect 19574 57692 19882 57712
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57616 19882 57636
rect 20444 57384 20496 57390
rect 20444 57326 20496 57332
rect 19574 56604 19882 56624
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56528 19882 56548
rect 19340 56296 19392 56302
rect 19340 56238 19392 56244
rect 19340 56160 19392 56166
rect 19340 56102 19392 56108
rect 17868 55208 17920 55214
rect 17868 55150 17920 55156
rect 19248 55208 19300 55214
rect 19248 55150 19300 55156
rect 19352 54874 19380 56102
rect 20456 55894 20484 57326
rect 22008 57316 22060 57322
rect 22008 57258 22060 57264
rect 22020 56370 22048 57258
rect 22560 56840 22612 56846
rect 22560 56782 22612 56788
rect 27252 56840 27304 56846
rect 27252 56782 27304 56788
rect 27896 56840 27948 56846
rect 27896 56782 27948 56788
rect 28264 56840 28316 56846
rect 28264 56782 28316 56788
rect 22376 56704 22428 56710
rect 22376 56646 22428 56652
rect 22388 56438 22416 56646
rect 22572 56506 22600 56782
rect 27160 56704 27212 56710
rect 27160 56646 27212 56652
rect 22560 56500 22612 56506
rect 22560 56442 22612 56448
rect 26976 56500 27028 56506
rect 26976 56442 27028 56448
rect 22376 56432 22428 56438
rect 22376 56374 22428 56380
rect 22008 56364 22060 56370
rect 22008 56306 22060 56312
rect 26148 56364 26200 56370
rect 26148 56306 26200 56312
rect 21824 56296 21876 56302
rect 21824 56238 21876 56244
rect 23020 56296 23072 56302
rect 23020 56238 23072 56244
rect 20444 55888 20496 55894
rect 20444 55830 20496 55836
rect 21836 55758 21864 56238
rect 23032 55826 23060 56238
rect 25596 56160 25648 56166
rect 25596 56102 25648 56108
rect 23020 55820 23072 55826
rect 23020 55762 23072 55768
rect 21824 55752 21876 55758
rect 21824 55694 21876 55700
rect 25044 55752 25096 55758
rect 25044 55694 25096 55700
rect 21272 55616 21324 55622
rect 21272 55558 21324 55564
rect 19574 55516 19882 55536
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55440 19882 55460
rect 21284 55282 21312 55558
rect 21836 55418 21864 55694
rect 22560 55616 22612 55622
rect 22560 55558 22612 55564
rect 21824 55412 21876 55418
rect 21824 55354 21876 55360
rect 22572 55350 22600 55558
rect 23664 55412 23716 55418
rect 23664 55354 23716 55360
rect 22560 55344 22612 55350
rect 22560 55286 22612 55292
rect 21272 55276 21324 55282
rect 21272 55218 21324 55224
rect 21916 55276 21968 55282
rect 21916 55218 21968 55224
rect 21088 55072 21140 55078
rect 21088 55014 21140 55020
rect 19340 54868 19392 54874
rect 19340 54810 19392 54816
rect 19156 54664 19208 54670
rect 19156 54606 19208 54612
rect 18696 50720 18748 50726
rect 18696 50662 18748 50668
rect 18708 50318 18736 50662
rect 18696 50312 18748 50318
rect 18696 50254 18748 50260
rect 19168 48822 19196 54606
rect 21100 54602 21128 55014
rect 21928 54670 21956 55218
rect 21916 54664 21968 54670
rect 21916 54606 21968 54612
rect 21088 54596 21140 54602
rect 21088 54538 21140 54544
rect 19984 54528 20036 54534
rect 19984 54470 20036 54476
rect 19574 54428 19882 54448
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54352 19882 54372
rect 19574 53340 19882 53360
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53264 19882 53284
rect 19574 52252 19882 52272
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52176 19882 52196
rect 19996 52018 20024 54470
rect 21928 53106 21956 54606
rect 22560 53576 22612 53582
rect 22560 53518 22612 53524
rect 22744 53576 22796 53582
rect 22744 53518 22796 53524
rect 22376 53440 22428 53446
rect 22376 53382 22428 53388
rect 21916 53100 21968 53106
rect 21916 53042 21968 53048
rect 22100 53100 22152 53106
rect 22100 53042 22152 53048
rect 21928 52494 21956 53042
rect 22112 52714 22140 53042
rect 22112 52686 22232 52714
rect 22100 52624 22152 52630
rect 22100 52566 22152 52572
rect 21916 52488 21968 52494
rect 21916 52430 21968 52436
rect 21928 52018 21956 52430
rect 22112 52086 22140 52566
rect 22100 52080 22152 52086
rect 22100 52022 22152 52028
rect 19984 52012 20036 52018
rect 19984 51954 20036 51960
rect 20076 52012 20128 52018
rect 20076 51954 20128 51960
rect 21916 52012 21968 52018
rect 21916 51954 21968 51960
rect 19340 51808 19392 51814
rect 19340 51750 19392 51756
rect 19352 51406 19380 51750
rect 19248 51400 19300 51406
rect 19248 51342 19300 51348
rect 19340 51400 19392 51406
rect 19340 51342 19392 51348
rect 19260 50386 19288 51342
rect 19574 51164 19882 51184
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51088 19882 51108
rect 19248 50380 19300 50386
rect 19248 50322 19300 50328
rect 19260 49434 19288 50322
rect 19574 50076 19882 50096
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50000 19882 50020
rect 19996 49978 20024 51954
rect 20088 50930 20116 51954
rect 22204 51610 22232 52686
rect 22192 51604 22244 51610
rect 22192 51546 22244 51552
rect 22388 51406 22416 53382
rect 22468 52420 22520 52426
rect 22468 52362 22520 52368
rect 22376 51400 22428 51406
rect 22376 51342 22428 51348
rect 20628 51264 20680 51270
rect 20628 51206 20680 51212
rect 20640 50998 20668 51206
rect 22480 51066 22508 52362
rect 22572 52154 22600 53518
rect 22652 52352 22704 52358
rect 22652 52294 22704 52300
rect 22560 52148 22612 52154
rect 22560 52090 22612 52096
rect 22664 51610 22692 52294
rect 22652 51604 22704 51610
rect 22652 51546 22704 51552
rect 22756 51406 22784 53518
rect 23676 53106 23704 55354
rect 25056 53650 25084 55694
rect 25412 55684 25464 55690
rect 25412 55626 25464 55632
rect 25424 55418 25452 55626
rect 25412 55412 25464 55418
rect 25412 55354 25464 55360
rect 25608 55282 25636 56102
rect 26160 55282 26188 56306
rect 26988 56302 27016 56442
rect 26976 56296 27028 56302
rect 26976 56238 27028 56244
rect 26332 55616 26384 55622
rect 26332 55558 26384 55564
rect 25596 55276 25648 55282
rect 25596 55218 25648 55224
rect 26148 55276 26200 55282
rect 26148 55218 26200 55224
rect 26056 55208 26108 55214
rect 26056 55150 26108 55156
rect 26068 54738 26096 55150
rect 26056 54732 26108 54738
rect 26056 54674 26108 54680
rect 26160 54194 26188 55218
rect 26344 54262 26372 55558
rect 26988 54602 27016 56238
rect 27172 55758 27200 56646
rect 27264 56506 27292 56782
rect 27252 56500 27304 56506
rect 27252 56442 27304 56448
rect 27908 56370 27936 56782
rect 28172 56704 28224 56710
rect 28172 56646 28224 56652
rect 28184 56438 28212 56646
rect 28172 56432 28224 56438
rect 28172 56374 28224 56380
rect 27896 56364 27948 56370
rect 27896 56306 27948 56312
rect 28276 56250 28304 56782
rect 28368 56302 28396 59200
rect 30196 56840 30248 56846
rect 30196 56782 30248 56788
rect 27620 56228 27672 56234
rect 27620 56170 27672 56176
rect 28184 56222 28304 56250
rect 28356 56296 28408 56302
rect 28356 56238 28408 56244
rect 27160 55752 27212 55758
rect 27160 55694 27212 55700
rect 27344 55344 27396 55350
rect 27396 55292 27568 55298
rect 27344 55286 27568 55292
rect 27356 55270 27568 55286
rect 27540 54754 27568 55270
rect 27632 55078 27660 56170
rect 28184 55894 28212 56222
rect 28172 55888 28224 55894
rect 28172 55830 28224 55836
rect 27620 55072 27672 55078
rect 27620 55014 27672 55020
rect 28080 55072 28132 55078
rect 28080 55014 28132 55020
rect 27632 54874 27660 55014
rect 27620 54868 27672 54874
rect 27620 54810 27672 54816
rect 27896 54868 27948 54874
rect 27896 54810 27948 54816
rect 27540 54726 27660 54754
rect 26976 54596 27028 54602
rect 26976 54538 27028 54544
rect 27436 54528 27488 54534
rect 27436 54470 27488 54476
rect 26332 54256 26384 54262
rect 26332 54198 26384 54204
rect 26148 54188 26200 54194
rect 26148 54130 26200 54136
rect 25044 53644 25096 53650
rect 25044 53586 25096 53592
rect 23664 53100 23716 53106
rect 23664 53042 23716 53048
rect 23204 52896 23256 52902
rect 23204 52838 23256 52844
rect 23480 52896 23532 52902
rect 23480 52838 23532 52844
rect 23112 52148 23164 52154
rect 23112 52090 23164 52096
rect 22744 51400 22796 51406
rect 22744 51342 22796 51348
rect 22468 51060 22520 51066
rect 22468 51002 22520 51008
rect 20260 50992 20312 50998
rect 20260 50934 20312 50940
rect 20628 50992 20680 50998
rect 20628 50934 20680 50940
rect 20076 50924 20128 50930
rect 20076 50866 20128 50872
rect 19432 49972 19484 49978
rect 19432 49914 19484 49920
rect 19984 49972 20036 49978
rect 19984 49914 20036 49920
rect 19248 49428 19300 49434
rect 19248 49370 19300 49376
rect 19260 49298 19288 49370
rect 19248 49292 19300 49298
rect 19248 49234 19300 49240
rect 19444 49162 19472 49914
rect 19432 49156 19484 49162
rect 19432 49098 19484 49104
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 19156 48816 19208 48822
rect 19156 48758 19208 48764
rect 19168 48074 19196 48758
rect 19708 48680 19760 48686
rect 19708 48622 19760 48628
rect 19720 48142 19748 48622
rect 19996 48550 20024 49914
rect 20088 49842 20116 50866
rect 20272 49910 20300 50934
rect 22756 50862 22784 51342
rect 23124 51338 23152 52090
rect 23216 52018 23244 52838
rect 23204 52012 23256 52018
rect 23204 51954 23256 51960
rect 23216 51474 23244 51954
rect 23204 51468 23256 51474
rect 23204 51410 23256 51416
rect 23112 51332 23164 51338
rect 23112 51274 23164 51280
rect 23216 50998 23244 51410
rect 23204 50992 23256 50998
rect 23204 50934 23256 50940
rect 23492 50930 23520 52838
rect 23676 52154 23704 53042
rect 25056 52562 25084 53586
rect 25412 53508 25464 53514
rect 25412 53450 25464 53456
rect 25424 53242 25452 53450
rect 26160 53258 26188 54130
rect 26240 53984 26292 53990
rect 26240 53926 26292 53932
rect 25412 53236 25464 53242
rect 25412 53178 25464 53184
rect 26068 53230 26188 53258
rect 25780 53168 25832 53174
rect 25780 53110 25832 53116
rect 25504 53100 25556 53106
rect 25504 53042 25556 53048
rect 25044 52556 25096 52562
rect 25044 52498 25096 52504
rect 23756 52352 23808 52358
rect 23756 52294 23808 52300
rect 23664 52148 23716 52154
rect 23664 52090 23716 52096
rect 23676 51610 23704 52090
rect 23768 51882 23796 52294
rect 25056 52018 25084 52498
rect 25044 52012 25096 52018
rect 25044 51954 25096 51960
rect 23756 51876 23808 51882
rect 23756 51818 23808 51824
rect 23664 51604 23716 51610
rect 23664 51546 23716 51552
rect 23768 51406 23796 51818
rect 24216 51808 24268 51814
rect 24216 51750 24268 51756
rect 23756 51400 23808 51406
rect 23756 51342 23808 51348
rect 23480 50924 23532 50930
rect 23480 50866 23532 50872
rect 22744 50856 22796 50862
rect 22744 50798 22796 50804
rect 23480 50788 23532 50794
rect 23480 50730 23532 50736
rect 22376 50720 22428 50726
rect 22376 50662 22428 50668
rect 22388 50318 22416 50662
rect 22376 50312 22428 50318
rect 22376 50254 22428 50260
rect 20628 50176 20680 50182
rect 20628 50118 20680 50124
rect 22192 50176 22244 50182
rect 22192 50118 22244 50124
rect 20640 49978 20668 50118
rect 20628 49972 20680 49978
rect 20628 49914 20680 49920
rect 20260 49904 20312 49910
rect 20260 49846 20312 49852
rect 20076 49836 20128 49842
rect 20076 49778 20128 49784
rect 20168 49768 20220 49774
rect 20168 49710 20220 49716
rect 20180 48822 20208 49710
rect 20272 48822 20300 49846
rect 20536 49836 20588 49842
rect 20536 49778 20588 49784
rect 20548 49450 20576 49778
rect 20640 49774 20668 49914
rect 20628 49768 20680 49774
rect 20628 49710 20680 49716
rect 22008 49768 22060 49774
rect 22008 49710 22060 49716
rect 20548 49422 20668 49450
rect 20640 49094 20668 49422
rect 21640 49224 21692 49230
rect 21640 49166 21692 49172
rect 20628 49088 20680 49094
rect 20628 49030 20680 49036
rect 20168 48816 20220 48822
rect 20168 48758 20220 48764
rect 20260 48816 20312 48822
rect 20260 48758 20312 48764
rect 20640 48686 20668 49030
rect 21652 48822 21680 49166
rect 21640 48816 21692 48822
rect 21640 48758 21692 48764
rect 20628 48680 20680 48686
rect 20628 48622 20680 48628
rect 19984 48544 20036 48550
rect 19984 48486 20036 48492
rect 21364 48544 21416 48550
rect 21364 48486 21416 48492
rect 19708 48136 19760 48142
rect 19708 48078 19760 48084
rect 19984 48136 20036 48142
rect 19984 48078 20036 48084
rect 19156 48068 19208 48074
rect 19156 48010 19208 48016
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 18788 47592 18840 47598
rect 18788 47534 18840 47540
rect 18800 46578 18828 47534
rect 19524 47456 19576 47462
rect 19524 47398 19576 47404
rect 19536 47122 19564 47398
rect 19524 47116 19576 47122
rect 19524 47058 19576 47064
rect 19996 47054 20024 48078
rect 20812 48000 20864 48006
rect 20812 47942 20864 47948
rect 20824 47666 20852 47942
rect 20812 47660 20864 47666
rect 20812 47602 20864 47608
rect 20168 47456 20220 47462
rect 20168 47398 20220 47404
rect 20076 47116 20128 47122
rect 20076 47058 20128 47064
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 19984 47048 20036 47054
rect 19984 46990 20036 46996
rect 18788 46572 18840 46578
rect 18788 46514 18840 46520
rect 18800 46034 18828 46514
rect 19352 46050 19380 46990
rect 19432 46980 19484 46986
rect 19432 46922 19484 46928
rect 18788 46028 18840 46034
rect 18788 45970 18840 45976
rect 19168 46022 19380 46050
rect 18800 45490 18828 45970
rect 19168 45966 19196 46022
rect 19156 45960 19208 45966
rect 19156 45902 19208 45908
rect 19340 45892 19392 45898
rect 19340 45834 19392 45840
rect 18788 45484 18840 45490
rect 18788 45426 18840 45432
rect 19352 45082 19380 45834
rect 19340 45076 19392 45082
rect 19340 45018 19392 45024
rect 19444 44878 19472 46922
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19984 46640 20036 46646
rect 19984 46582 20036 46588
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19996 44538 20024 46582
rect 19984 44532 20036 44538
rect 19984 44474 20036 44480
rect 20088 44402 20116 47058
rect 20180 45354 20208 47398
rect 21376 47054 21404 48486
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 21364 47048 21416 47054
rect 21364 46990 21416 46996
rect 20260 46096 20312 46102
rect 20260 46038 20312 46044
rect 20272 45490 20300 46038
rect 20260 45484 20312 45490
rect 20260 45426 20312 45432
rect 20168 45348 20220 45354
rect 20168 45290 20220 45296
rect 20180 45082 20208 45290
rect 20364 45286 20392 46990
rect 20628 46980 20680 46986
rect 20628 46922 20680 46928
rect 20444 46368 20496 46374
rect 20444 46310 20496 46316
rect 20456 45626 20484 46310
rect 20536 46164 20588 46170
rect 20536 46106 20588 46112
rect 20444 45620 20496 45626
rect 20444 45562 20496 45568
rect 20352 45280 20404 45286
rect 20352 45222 20404 45228
rect 20168 45076 20220 45082
rect 20168 45018 20220 45024
rect 20364 44826 20392 45222
rect 20456 44946 20484 45562
rect 20548 45490 20576 46106
rect 20536 45484 20588 45490
rect 20536 45426 20588 45432
rect 20444 44940 20496 44946
rect 20444 44882 20496 44888
rect 20548 44878 20576 45426
rect 20640 45082 20668 46922
rect 22020 46578 22048 49710
rect 22204 49230 22232 50118
rect 23492 49858 23520 50730
rect 24032 49904 24084 49910
rect 23492 49842 23704 49858
rect 24032 49846 24084 49852
rect 23480 49836 23704 49842
rect 23532 49830 23704 49836
rect 23480 49778 23532 49784
rect 23572 49768 23624 49774
rect 23572 49710 23624 49716
rect 23480 49700 23532 49706
rect 23480 49642 23532 49648
rect 22376 49632 22428 49638
rect 22376 49574 22428 49580
rect 22192 49224 22244 49230
rect 22192 49166 22244 49172
rect 22388 48754 22416 49574
rect 23492 48890 23520 49642
rect 23584 49434 23612 49710
rect 23572 49428 23624 49434
rect 23572 49370 23624 49376
rect 23676 49230 23704 49830
rect 23848 49768 23900 49774
rect 23848 49710 23900 49716
rect 23664 49224 23716 49230
rect 23664 49166 23716 49172
rect 23756 49156 23808 49162
rect 23756 49098 23808 49104
rect 23480 48884 23532 48890
rect 23480 48826 23532 48832
rect 22376 48748 22428 48754
rect 22376 48690 22428 48696
rect 23768 48346 23796 49098
rect 23756 48340 23808 48346
rect 23756 48282 23808 48288
rect 23860 48142 23888 49710
rect 24044 49094 24072 49846
rect 24124 49836 24176 49842
rect 24124 49778 24176 49784
rect 24136 49298 24164 49778
rect 24124 49292 24176 49298
rect 24124 49234 24176 49240
rect 24032 49088 24084 49094
rect 24032 49030 24084 49036
rect 24044 48754 24072 49030
rect 24032 48748 24084 48754
rect 24032 48690 24084 48696
rect 24136 48550 24164 49234
rect 24124 48544 24176 48550
rect 24124 48486 24176 48492
rect 23848 48136 23900 48142
rect 23848 48078 23900 48084
rect 24228 47666 24256 51750
rect 24584 51264 24636 51270
rect 24584 51206 24636 51212
rect 24400 49836 24452 49842
rect 24400 49778 24452 49784
rect 24308 48884 24360 48890
rect 24308 48826 24360 48832
rect 24320 48754 24348 48826
rect 24308 48748 24360 48754
rect 24308 48690 24360 48696
rect 24412 48686 24440 49778
rect 24400 48680 24452 48686
rect 24400 48622 24452 48628
rect 24400 48544 24452 48550
rect 24400 48486 24452 48492
rect 24412 48142 24440 48486
rect 24596 48142 24624 51206
rect 25056 50522 25084 51954
rect 25516 51338 25544 53042
rect 25792 51406 25820 53110
rect 25780 51400 25832 51406
rect 25780 51342 25832 51348
rect 25504 51332 25556 51338
rect 25504 51274 25556 51280
rect 25516 50930 25544 51274
rect 25504 50924 25556 50930
rect 25504 50866 25556 50872
rect 25596 50856 25648 50862
rect 25596 50798 25648 50804
rect 25044 50516 25096 50522
rect 25044 50458 25096 50464
rect 24676 49768 24728 49774
rect 24676 49710 24728 49716
rect 24400 48136 24452 48142
rect 24400 48078 24452 48084
rect 24584 48136 24636 48142
rect 24584 48078 24636 48084
rect 24688 47802 24716 49710
rect 25056 49230 25084 50458
rect 25608 50318 25636 50798
rect 25792 50726 25820 51342
rect 25780 50720 25832 50726
rect 25780 50662 25832 50668
rect 25596 50312 25648 50318
rect 25596 50254 25648 50260
rect 25608 49774 25636 50254
rect 25792 49774 25820 50662
rect 26068 50386 26096 53230
rect 26252 53122 26280 53926
rect 26344 53718 26372 54198
rect 27448 53786 27476 54470
rect 27436 53780 27488 53786
rect 27436 53722 27488 53728
rect 26332 53712 26384 53718
rect 26332 53654 26384 53660
rect 27252 53712 27304 53718
rect 27252 53654 27304 53660
rect 26792 53576 26844 53582
rect 26792 53518 26844 53524
rect 26160 53106 26280 53122
rect 26148 53100 26280 53106
rect 26200 53094 26280 53100
rect 26148 53042 26200 53048
rect 26804 53038 26832 53518
rect 26884 53508 26936 53514
rect 26884 53450 26936 53456
rect 26896 53106 26924 53450
rect 27160 53440 27212 53446
rect 27160 53382 27212 53388
rect 26884 53100 26936 53106
rect 26884 53042 26936 53048
rect 26792 53032 26844 53038
rect 26792 52974 26844 52980
rect 26424 52896 26476 52902
rect 26424 52838 26476 52844
rect 26436 52018 26464 52838
rect 26804 52154 26832 52974
rect 26896 52630 26924 53042
rect 27172 52970 27200 53382
rect 27264 53106 27292 53654
rect 27436 53576 27488 53582
rect 27436 53518 27488 53524
rect 27448 53242 27476 53518
rect 27436 53236 27488 53242
rect 27436 53178 27488 53184
rect 27252 53100 27304 53106
rect 27252 53042 27304 53048
rect 27344 53100 27396 53106
rect 27344 53042 27396 53048
rect 27160 52964 27212 52970
rect 27160 52906 27212 52912
rect 27068 52896 27120 52902
rect 27068 52838 27120 52844
rect 26884 52624 26936 52630
rect 26884 52566 26936 52572
rect 26792 52148 26844 52154
rect 26792 52090 26844 52096
rect 26424 52012 26476 52018
rect 26424 51954 26476 51960
rect 26896 51474 26924 52566
rect 26976 52488 27028 52494
rect 26976 52430 27028 52436
rect 26988 52154 27016 52430
rect 26976 52148 27028 52154
rect 26976 52090 27028 52096
rect 27080 52086 27108 52838
rect 27068 52080 27120 52086
rect 27068 52022 27120 52028
rect 27356 51610 27384 53042
rect 27344 51604 27396 51610
rect 27344 51546 27396 51552
rect 26884 51468 26936 51474
rect 26884 51410 26936 51416
rect 26056 50380 26108 50386
rect 26056 50322 26108 50328
rect 25964 50244 26016 50250
rect 25964 50186 26016 50192
rect 25596 49768 25648 49774
rect 25596 49710 25648 49716
rect 25780 49768 25832 49774
rect 25780 49710 25832 49716
rect 25044 49224 25096 49230
rect 25044 49166 25096 49172
rect 25056 48754 25084 49166
rect 25044 48748 25096 48754
rect 25044 48690 25096 48696
rect 25608 48210 25636 49710
rect 25596 48204 25648 48210
rect 25596 48146 25648 48152
rect 24768 48000 24820 48006
rect 24768 47942 24820 47948
rect 24676 47796 24728 47802
rect 24676 47738 24728 47744
rect 24780 47734 24808 47942
rect 24768 47728 24820 47734
rect 24768 47670 24820 47676
rect 24216 47660 24268 47666
rect 24216 47602 24268 47608
rect 24676 47592 24728 47598
rect 24676 47534 24728 47540
rect 24492 47456 24544 47462
rect 24492 47398 24544 47404
rect 24504 47054 24532 47398
rect 24032 47048 24084 47054
rect 24032 46990 24084 46996
rect 24400 47048 24452 47054
rect 24400 46990 24452 46996
rect 24492 47048 24544 47054
rect 24492 46990 24544 46996
rect 22284 46980 22336 46986
rect 22284 46922 22336 46928
rect 22296 46646 22324 46922
rect 22652 46912 22704 46918
rect 22652 46854 22704 46860
rect 22284 46640 22336 46646
rect 22284 46582 22336 46588
rect 22664 46578 22692 46854
rect 24044 46714 24072 46990
rect 24032 46708 24084 46714
rect 24032 46650 24084 46656
rect 22008 46572 22060 46578
rect 22008 46514 22060 46520
rect 22100 46572 22152 46578
rect 22100 46514 22152 46520
rect 22652 46572 22704 46578
rect 22652 46514 22704 46520
rect 21824 46368 21876 46374
rect 21824 46310 21876 46316
rect 21836 45898 21864 46310
rect 21824 45892 21876 45898
rect 21824 45834 21876 45840
rect 22112 45490 22140 46514
rect 22376 45960 22428 45966
rect 22376 45902 22428 45908
rect 22100 45484 22152 45490
rect 22100 45426 22152 45432
rect 22388 45422 22416 45902
rect 22664 45558 22692 46514
rect 23664 46504 23716 46510
rect 23664 46446 23716 46452
rect 23112 46368 23164 46374
rect 23112 46310 23164 46316
rect 23124 45966 23152 46310
rect 23676 46102 23704 46446
rect 23664 46096 23716 46102
rect 23664 46038 23716 46044
rect 24216 46096 24268 46102
rect 24216 46038 24268 46044
rect 23112 45960 23164 45966
rect 23112 45902 23164 45908
rect 22652 45552 22704 45558
rect 22652 45494 22704 45500
rect 24228 45422 24256 46038
rect 24412 46034 24440 46990
rect 24400 46028 24452 46034
rect 24400 45970 24452 45976
rect 24688 45898 24716 47534
rect 25976 47462 26004 50186
rect 26068 49298 26096 50322
rect 27632 49910 27660 54726
rect 27908 54194 27936 54810
rect 28092 54602 28120 55014
rect 28080 54596 28132 54602
rect 28080 54538 28132 54544
rect 27896 54188 27948 54194
rect 27896 54130 27948 54136
rect 28184 53174 28212 55830
rect 30208 55826 30236 56782
rect 30300 55826 30328 59200
rect 31588 57882 31616 59200
rect 31588 57854 31800 57882
rect 31300 57248 31352 57254
rect 31300 57190 31352 57196
rect 31312 56846 31340 57190
rect 30656 56840 30708 56846
rect 30656 56782 30708 56788
rect 31300 56840 31352 56846
rect 31300 56782 31352 56788
rect 30668 56438 30696 56782
rect 31772 56778 31800 57854
rect 32128 57248 32180 57254
rect 32128 57190 32180 57196
rect 31760 56772 31812 56778
rect 31760 56714 31812 56720
rect 30656 56432 30708 56438
rect 30656 56374 30708 56380
rect 31484 56432 31536 56438
rect 31484 56374 31536 56380
rect 30932 56160 30984 56166
rect 30932 56102 30984 56108
rect 30196 55820 30248 55826
rect 30196 55762 30248 55768
rect 30288 55820 30340 55826
rect 30288 55762 30340 55768
rect 30944 55690 30972 56102
rect 30932 55684 30984 55690
rect 30932 55626 30984 55632
rect 28448 55616 28500 55622
rect 28448 55558 28500 55564
rect 28460 54874 28488 55558
rect 28540 55344 28592 55350
rect 28540 55286 28592 55292
rect 28552 55214 28580 55286
rect 29276 55276 29328 55282
rect 29276 55218 29328 55224
rect 28540 55208 28592 55214
rect 28540 55150 28592 55156
rect 29288 55146 29316 55218
rect 29552 55208 29604 55214
rect 29552 55150 29604 55156
rect 29276 55140 29328 55146
rect 29276 55082 29328 55088
rect 28448 54868 28500 54874
rect 28448 54810 28500 54816
rect 29000 54732 29052 54738
rect 29000 54674 29052 54680
rect 29012 54534 29040 54674
rect 29564 54670 29592 55150
rect 29552 54664 29604 54670
rect 29552 54606 29604 54612
rect 28448 54528 28500 54534
rect 28448 54470 28500 54476
rect 28724 54528 28776 54534
rect 28724 54470 28776 54476
rect 29000 54528 29052 54534
rect 29000 54470 29052 54476
rect 28460 54194 28488 54470
rect 28448 54188 28500 54194
rect 28448 54130 28500 54136
rect 28736 53582 28764 54470
rect 29012 54126 29040 54470
rect 29184 54256 29236 54262
rect 29184 54198 29236 54204
rect 29000 54120 29052 54126
rect 29000 54062 29052 54068
rect 29092 54120 29144 54126
rect 29092 54062 29144 54068
rect 29104 53786 29132 54062
rect 29092 53780 29144 53786
rect 29092 53722 29144 53728
rect 28724 53576 28776 53582
rect 28724 53518 28776 53524
rect 29000 53576 29052 53582
rect 29000 53518 29052 53524
rect 28448 53508 28500 53514
rect 28448 53450 28500 53456
rect 28172 53168 28224 53174
rect 28172 53110 28224 53116
rect 28460 51074 28488 53450
rect 29012 52494 29040 53518
rect 29000 52488 29052 52494
rect 29000 52430 29052 52436
rect 29000 52012 29052 52018
rect 29000 51954 29052 51960
rect 28816 51264 28868 51270
rect 28816 51206 28868 51212
rect 28460 51046 28580 51074
rect 28264 50924 28316 50930
rect 28264 50866 28316 50872
rect 28276 50318 28304 50866
rect 28264 50312 28316 50318
rect 28264 50254 28316 50260
rect 27620 49904 27672 49910
rect 27620 49846 27672 49852
rect 28276 49842 28304 50254
rect 28264 49836 28316 49842
rect 28264 49778 28316 49784
rect 26056 49292 26108 49298
rect 26056 49234 26108 49240
rect 28276 49230 28304 49778
rect 28264 49224 28316 49230
rect 28264 49166 28316 49172
rect 27896 49156 27948 49162
rect 27896 49098 27948 49104
rect 27160 49088 27212 49094
rect 27160 49030 27212 49036
rect 27172 48754 27200 49030
rect 27908 48890 27936 49098
rect 27896 48884 27948 48890
rect 27896 48826 27948 48832
rect 27160 48748 27212 48754
rect 27160 48690 27212 48696
rect 28080 48748 28132 48754
rect 28080 48690 28132 48696
rect 26976 48272 27028 48278
rect 26976 48214 27028 48220
rect 26148 48136 26200 48142
rect 26148 48078 26200 48084
rect 26160 47666 26188 48078
rect 26056 47660 26108 47666
rect 26056 47602 26108 47608
rect 26148 47660 26200 47666
rect 26148 47602 26200 47608
rect 25964 47456 26016 47462
rect 25964 47398 26016 47404
rect 25780 46912 25832 46918
rect 25780 46854 25832 46860
rect 24860 46708 24912 46714
rect 24860 46650 24912 46656
rect 24872 46578 24900 46650
rect 24860 46572 24912 46578
rect 24860 46514 24912 46520
rect 25792 46510 25820 46854
rect 25976 46646 26004 47398
rect 25964 46640 26016 46646
rect 25964 46582 26016 46588
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 25780 46504 25832 46510
rect 25780 46446 25832 46452
rect 25964 46504 26016 46510
rect 25964 46446 26016 46452
rect 24952 46368 25004 46374
rect 24952 46310 25004 46316
rect 24964 45966 24992 46310
rect 24952 45960 25004 45966
rect 24952 45902 25004 45908
rect 24676 45892 24728 45898
rect 24676 45834 24728 45840
rect 25148 45558 25176 46446
rect 25596 45824 25648 45830
rect 25596 45766 25648 45772
rect 25608 45558 25636 45766
rect 25136 45552 25188 45558
rect 25136 45494 25188 45500
rect 25596 45552 25648 45558
rect 25596 45494 25648 45500
rect 22376 45416 22428 45422
rect 22376 45358 22428 45364
rect 24216 45416 24268 45422
rect 24216 45358 24268 45364
rect 20628 45076 20680 45082
rect 20628 45018 20680 45024
rect 20272 44810 20392 44826
rect 20536 44872 20588 44878
rect 20536 44814 20588 44820
rect 20260 44804 20392 44810
rect 20312 44798 20392 44804
rect 20260 44746 20312 44752
rect 20076 44396 20128 44402
rect 20076 44338 20128 44344
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 21456 42900 21508 42906
rect 21456 42842 21508 42848
rect 20628 42764 20680 42770
rect 20628 42706 20680 42712
rect 20260 42696 20312 42702
rect 20260 42638 20312 42644
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 20272 42362 20300 42638
rect 20260 42356 20312 42362
rect 20260 42298 20312 42304
rect 20168 42220 20220 42226
rect 20168 42162 20220 42168
rect 20180 41818 20208 42162
rect 20640 42158 20668 42706
rect 21180 42696 21232 42702
rect 21180 42638 21232 42644
rect 21192 42294 21220 42638
rect 21272 42628 21324 42634
rect 21272 42570 21324 42576
rect 21180 42288 21232 42294
rect 21180 42230 21232 42236
rect 20628 42152 20680 42158
rect 20628 42094 20680 42100
rect 21284 41818 21312 42570
rect 20168 41812 20220 41818
rect 20168 41754 20220 41760
rect 20996 41812 21048 41818
rect 20996 41754 21048 41760
rect 21272 41812 21324 41818
rect 21272 41754 21324 41760
rect 20442 41712 20498 41721
rect 20442 41647 20498 41656
rect 20456 41614 20484 41647
rect 19984 41608 20036 41614
rect 19984 41550 20036 41556
rect 20444 41608 20496 41614
rect 20812 41608 20864 41614
rect 20444 41550 20496 41556
rect 20810 41576 20812 41585
rect 20864 41576 20866 41585
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19996 41002 20024 41550
rect 20810 41511 20866 41520
rect 21008 41070 21036 41754
rect 21180 41676 21232 41682
rect 21180 41618 21232 41624
rect 21088 41472 21140 41478
rect 21088 41414 21140 41420
rect 20536 41064 20588 41070
rect 20536 41006 20588 41012
rect 20996 41064 21048 41070
rect 20996 41006 21048 41012
rect 19984 40996 20036 41002
rect 19984 40938 20036 40944
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 20548 40118 20576 41006
rect 21100 40730 21128 41414
rect 21088 40724 21140 40730
rect 21088 40666 21140 40672
rect 20536 40112 20588 40118
rect 20536 40054 20588 40060
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19524 38752 19576 38758
rect 19524 38694 19576 38700
rect 19536 38282 19564 38694
rect 19524 38276 19576 38282
rect 19524 38218 19576 38224
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 20548 37806 20576 40054
rect 20904 39432 20956 39438
rect 20904 39374 20956 39380
rect 20812 38752 20864 38758
rect 20812 38694 20864 38700
rect 20628 38344 20680 38350
rect 20628 38286 20680 38292
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20364 37262 20392 37606
rect 20640 37262 20668 38286
rect 20720 38208 20772 38214
rect 20720 38150 20772 38156
rect 20732 37874 20760 38150
rect 20720 37868 20772 37874
rect 20720 37810 20772 37816
rect 20824 37330 20852 38694
rect 20916 37466 20944 39374
rect 21088 39296 21140 39302
rect 21088 39238 21140 39244
rect 21100 38962 21128 39238
rect 21088 38956 21140 38962
rect 21088 38898 21140 38904
rect 21192 38894 21220 41618
rect 21468 41546 21496 42842
rect 22388 42294 22416 45358
rect 25148 45354 25176 45494
rect 25136 45348 25188 45354
rect 25136 45290 25188 45296
rect 24676 45280 24728 45286
rect 24676 45222 24728 45228
rect 24768 45280 24820 45286
rect 24768 45222 24820 45228
rect 24688 44878 24716 45222
rect 24780 44878 24808 45222
rect 24860 45076 24912 45082
rect 24860 45018 24912 45024
rect 24676 44872 24728 44878
rect 24676 44814 24728 44820
rect 24768 44872 24820 44878
rect 24768 44814 24820 44820
rect 24216 44736 24268 44742
rect 24216 44678 24268 44684
rect 24228 43382 24256 44678
rect 24688 44266 24716 44814
rect 24780 44538 24808 44814
rect 24768 44532 24820 44538
rect 24768 44474 24820 44480
rect 24872 44402 24900 45018
rect 25608 44878 25636 45494
rect 25688 45484 25740 45490
rect 25688 45426 25740 45432
rect 25700 44878 25728 45426
rect 25976 44962 26004 46446
rect 26068 46170 26096 47602
rect 26160 47054 26188 47602
rect 26148 47048 26200 47054
rect 26148 46990 26200 46996
rect 26160 46714 26188 46990
rect 26988 46918 27016 48214
rect 28092 48210 28120 48690
rect 28080 48204 28132 48210
rect 28080 48146 28132 48152
rect 27620 48136 27672 48142
rect 27620 48078 27672 48084
rect 27632 47666 27660 48078
rect 27620 47660 27672 47666
rect 27672 47620 27752 47648
rect 27620 47602 27672 47608
rect 27620 47456 27672 47462
rect 27620 47398 27672 47404
rect 27632 47122 27660 47398
rect 27620 47116 27672 47122
rect 27620 47058 27672 47064
rect 27160 47048 27212 47054
rect 27160 46990 27212 46996
rect 26976 46912 27028 46918
rect 26976 46854 27028 46860
rect 26148 46708 26200 46714
rect 26148 46650 26200 46656
rect 26424 46436 26476 46442
rect 26424 46378 26476 46384
rect 26056 46164 26108 46170
rect 26056 46106 26108 46112
rect 26056 45280 26108 45286
rect 26056 45222 26108 45228
rect 26068 45082 26096 45222
rect 26056 45076 26108 45082
rect 26056 45018 26108 45024
rect 25976 44934 26096 44962
rect 25044 44872 25096 44878
rect 25044 44814 25096 44820
rect 25596 44872 25648 44878
rect 25596 44814 25648 44820
rect 25688 44872 25740 44878
rect 25688 44814 25740 44820
rect 25056 44402 25084 44814
rect 24860 44396 24912 44402
rect 24860 44338 24912 44344
rect 25044 44396 25096 44402
rect 25044 44338 25096 44344
rect 24676 44260 24728 44266
rect 24676 44202 24728 44208
rect 24400 44192 24452 44198
rect 24400 44134 24452 44140
rect 24216 43376 24268 43382
rect 24216 43318 24268 43324
rect 23296 43308 23348 43314
rect 23296 43250 23348 43256
rect 22560 43104 22612 43110
rect 22560 43046 22612 43052
rect 22376 42288 22428 42294
rect 22376 42230 22428 42236
rect 22008 42220 22060 42226
rect 22008 42162 22060 42168
rect 22020 41818 22048 42162
rect 22284 42016 22336 42022
rect 22284 41958 22336 41964
rect 22008 41812 22060 41818
rect 22008 41754 22060 41760
rect 21732 41608 21784 41614
rect 21916 41608 21968 41614
rect 21732 41550 21784 41556
rect 21914 41576 21916 41585
rect 22192 41608 22244 41614
rect 21968 41576 21970 41585
rect 21456 41540 21508 41546
rect 21456 41482 21508 41488
rect 21744 40730 21772 41550
rect 22192 41550 22244 41556
rect 21914 41511 21970 41520
rect 21824 41472 21876 41478
rect 21824 41414 21876 41420
rect 21836 40730 21864 41414
rect 22204 41274 22232 41550
rect 22192 41268 22244 41274
rect 22192 41210 22244 41216
rect 21732 40724 21784 40730
rect 21732 40666 21784 40672
rect 21824 40724 21876 40730
rect 21824 40666 21876 40672
rect 21916 40656 21968 40662
rect 21916 40598 21968 40604
rect 21928 40526 21956 40598
rect 21916 40520 21968 40526
rect 21916 40462 21968 40468
rect 21928 39506 21956 40462
rect 22204 40458 22232 41210
rect 22296 40594 22324 41958
rect 22572 41721 22600 43046
rect 23308 42838 23336 43250
rect 23480 43172 23532 43178
rect 23480 43114 23532 43120
rect 23388 43104 23440 43110
rect 23388 43046 23440 43052
rect 23400 42906 23428 43046
rect 23388 42900 23440 42906
rect 23388 42842 23440 42848
rect 22744 42832 22796 42838
rect 22744 42774 22796 42780
rect 23296 42832 23348 42838
rect 23296 42774 23348 42780
rect 22558 41712 22614 41721
rect 22376 41676 22428 41682
rect 22558 41647 22614 41656
rect 22376 41618 22428 41624
rect 22284 40588 22336 40594
rect 22284 40530 22336 40536
rect 22192 40452 22244 40458
rect 22192 40394 22244 40400
rect 22284 40384 22336 40390
rect 22284 40326 22336 40332
rect 22296 40118 22324 40326
rect 22284 40112 22336 40118
rect 22284 40054 22336 40060
rect 22192 40044 22244 40050
rect 22192 39986 22244 39992
rect 21916 39500 21968 39506
rect 21916 39442 21968 39448
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 21180 38888 21232 38894
rect 21180 38830 21232 38836
rect 20996 38820 21048 38826
rect 20996 38762 21048 38768
rect 21008 37670 21036 38762
rect 21192 38554 21220 38830
rect 21180 38548 21232 38554
rect 21180 38490 21232 38496
rect 22112 38214 22140 38898
rect 22204 38758 22232 39986
rect 22388 38962 22416 41618
rect 22376 38956 22428 38962
rect 22376 38898 22428 38904
rect 22284 38888 22336 38894
rect 22284 38830 22336 38836
rect 22192 38752 22244 38758
rect 22192 38694 22244 38700
rect 21640 38208 21692 38214
rect 21640 38150 21692 38156
rect 22100 38208 22152 38214
rect 22100 38150 22152 38156
rect 20996 37664 21048 37670
rect 20996 37606 21048 37612
rect 20904 37460 20956 37466
rect 20904 37402 20956 37408
rect 20812 37324 20864 37330
rect 20812 37266 20864 37272
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 21652 37194 21680 38150
rect 21640 37188 21692 37194
rect 21640 37130 21692 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 22204 36718 22232 38694
rect 22296 38486 22324 38830
rect 22284 38480 22336 38486
rect 22284 38422 22336 38428
rect 22388 38350 22416 38898
rect 22376 38344 22428 38350
rect 22376 38286 22428 38292
rect 22468 38276 22520 38282
rect 22468 38218 22520 38224
rect 22480 38010 22508 38218
rect 22468 38004 22520 38010
rect 22468 37946 22520 37952
rect 22376 37800 22428 37806
rect 22376 37742 22428 37748
rect 22388 37262 22416 37742
rect 22376 37256 22428 37262
rect 22376 37198 22428 37204
rect 22388 37126 22416 37198
rect 22376 37120 22428 37126
rect 22376 37062 22428 37068
rect 22388 36786 22416 37062
rect 22572 36854 22600 41647
rect 22756 41546 22784 42774
rect 23388 42764 23440 42770
rect 23388 42706 23440 42712
rect 22836 42696 22888 42702
rect 22836 42638 22888 42644
rect 22848 41614 22876 42638
rect 23400 42294 23428 42706
rect 23492 42702 23520 43114
rect 23664 42832 23716 42838
rect 23664 42774 23716 42780
rect 23480 42696 23532 42702
rect 23480 42638 23532 42644
rect 23492 42362 23520 42638
rect 23480 42356 23532 42362
rect 23480 42298 23532 42304
rect 23388 42288 23440 42294
rect 23388 42230 23440 42236
rect 22836 41608 22888 41614
rect 22836 41550 22888 41556
rect 22744 41540 22796 41546
rect 22744 41482 22796 41488
rect 22756 41206 22784 41482
rect 22744 41200 22796 41206
rect 22744 41142 22796 41148
rect 22652 40656 22704 40662
rect 22652 40598 22704 40604
rect 22664 38962 22692 40598
rect 22744 40452 22796 40458
rect 22744 40394 22796 40400
rect 22756 39438 22784 40394
rect 22848 40050 22876 41550
rect 23676 41070 23704 42774
rect 23756 42696 23808 42702
rect 23756 42638 23808 42644
rect 23664 41064 23716 41070
rect 23664 41006 23716 41012
rect 23664 40588 23716 40594
rect 23664 40530 23716 40536
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 23676 39982 23704 40530
rect 23768 40458 23796 42638
rect 23940 42220 23992 42226
rect 23940 42162 23992 42168
rect 23952 41818 23980 42162
rect 23940 41812 23992 41818
rect 23940 41754 23992 41760
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 24136 41138 24164 41550
rect 24228 41414 24256 43318
rect 24412 43246 24440 44134
rect 26068 43314 26096 44934
rect 26240 43376 26292 43382
rect 26240 43318 26292 43324
rect 25228 43308 25280 43314
rect 25228 43250 25280 43256
rect 26056 43308 26108 43314
rect 26056 43250 26108 43256
rect 24400 43240 24452 43246
rect 24400 43182 24452 43188
rect 24412 42922 24440 43182
rect 24492 43172 24544 43178
rect 24492 43114 24544 43120
rect 24320 42894 24440 42922
rect 24320 42702 24348 42894
rect 24504 42702 24532 43114
rect 24676 43104 24728 43110
rect 24676 43046 24728 43052
rect 24688 42702 24716 43046
rect 24952 42832 25004 42838
rect 24952 42774 25004 42780
rect 24308 42696 24360 42702
rect 24308 42638 24360 42644
rect 24492 42696 24544 42702
rect 24492 42638 24544 42644
rect 24676 42696 24728 42702
rect 24676 42638 24728 42644
rect 24492 42560 24544 42566
rect 24492 42502 24544 42508
rect 24228 41386 24440 41414
rect 23940 41132 23992 41138
rect 23940 41074 23992 41080
rect 24124 41132 24176 41138
rect 24124 41074 24176 41080
rect 23756 40452 23808 40458
rect 23756 40394 23808 40400
rect 23952 40186 23980 41074
rect 23940 40180 23992 40186
rect 23940 40122 23992 40128
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23940 39568 23992 39574
rect 23940 39510 23992 39516
rect 22744 39432 22796 39438
rect 22744 39374 22796 39380
rect 23848 39364 23900 39370
rect 23848 39306 23900 39312
rect 23388 39092 23440 39098
rect 23388 39034 23440 39040
rect 22836 39024 22888 39030
rect 22836 38966 22888 38972
rect 22652 38956 22704 38962
rect 22652 38898 22704 38904
rect 22664 38350 22692 38898
rect 22652 38344 22704 38350
rect 22652 38286 22704 38292
rect 22652 38208 22704 38214
rect 22652 38150 22704 38156
rect 22664 38010 22692 38150
rect 22652 38004 22704 38010
rect 22652 37946 22704 37952
rect 22664 37806 22692 37946
rect 22652 37800 22704 37806
rect 22652 37742 22704 37748
rect 22848 37670 22876 38966
rect 23400 38962 23428 39034
rect 23860 38962 23888 39306
rect 23388 38956 23440 38962
rect 23388 38898 23440 38904
rect 23848 38956 23900 38962
rect 23848 38898 23900 38904
rect 23204 38820 23256 38826
rect 23204 38762 23256 38768
rect 22928 38752 22980 38758
rect 22928 38694 22980 38700
rect 22940 38350 22968 38694
rect 23216 38350 23244 38762
rect 22928 38344 22980 38350
rect 22928 38286 22980 38292
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 22928 37800 22980 37806
rect 22928 37742 22980 37748
rect 22836 37664 22888 37670
rect 22836 37606 22888 37612
rect 22560 36848 22612 36854
rect 22560 36790 22612 36796
rect 22848 36786 22876 37606
rect 22940 36786 22968 37742
rect 22376 36780 22428 36786
rect 22376 36722 22428 36728
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 22928 36780 22980 36786
rect 22928 36722 22980 36728
rect 22192 36712 22244 36718
rect 22192 36654 22244 36660
rect 23216 36650 23244 38286
rect 23400 37466 23428 38898
rect 23860 38826 23888 38898
rect 23848 38820 23900 38826
rect 23848 38762 23900 38768
rect 23952 38758 23980 39510
rect 24136 39506 24164 41074
rect 24308 40520 24360 40526
rect 24308 40462 24360 40468
rect 24320 40118 24348 40462
rect 24308 40112 24360 40118
rect 24308 40054 24360 40060
rect 24320 39642 24348 40054
rect 24308 39636 24360 39642
rect 24308 39578 24360 39584
rect 24124 39500 24176 39506
rect 24124 39442 24176 39448
rect 24412 38894 24440 41386
rect 24504 40594 24532 42502
rect 24584 42016 24636 42022
rect 24584 41958 24636 41964
rect 24596 41478 24624 41958
rect 24964 41818 24992 42774
rect 25240 42362 25268 43250
rect 25964 43104 26016 43110
rect 25964 43046 26016 43052
rect 25780 42628 25832 42634
rect 25780 42570 25832 42576
rect 25792 42362 25820 42570
rect 25228 42356 25280 42362
rect 25228 42298 25280 42304
rect 25780 42356 25832 42362
rect 25780 42298 25832 42304
rect 24952 41812 25004 41818
rect 24952 41754 25004 41760
rect 25044 41676 25096 41682
rect 25044 41618 25096 41624
rect 24768 41540 24820 41546
rect 24768 41482 24820 41488
rect 24584 41472 24636 41478
rect 24584 41414 24636 41420
rect 24596 41138 24624 41414
rect 24584 41132 24636 41138
rect 24584 41074 24636 41080
rect 24780 41002 24808 41482
rect 25056 41478 25084 41618
rect 25240 41614 25268 42298
rect 25976 42226 26004 43046
rect 25964 42220 26016 42226
rect 25964 42162 26016 42168
rect 25228 41608 25280 41614
rect 25228 41550 25280 41556
rect 25044 41472 25096 41478
rect 25044 41414 25096 41420
rect 24860 41268 24912 41274
rect 24860 41210 24912 41216
rect 24768 40996 24820 41002
rect 24768 40938 24820 40944
rect 24676 40928 24728 40934
rect 24676 40870 24728 40876
rect 24492 40588 24544 40594
rect 24492 40530 24544 40536
rect 24492 40044 24544 40050
rect 24492 39986 24544 39992
rect 24504 39642 24532 39986
rect 24492 39636 24544 39642
rect 24492 39578 24544 39584
rect 24584 39636 24636 39642
rect 24584 39578 24636 39584
rect 24596 39438 24624 39578
rect 24584 39432 24636 39438
rect 24584 39374 24636 39380
rect 24688 38894 24716 40870
rect 24872 39438 24900 41210
rect 24952 41064 25004 41070
rect 24952 41006 25004 41012
rect 24860 39432 24912 39438
rect 24860 39374 24912 39380
rect 24400 38888 24452 38894
rect 24400 38830 24452 38836
rect 24676 38888 24728 38894
rect 24676 38830 24728 38836
rect 23940 38752 23992 38758
rect 23940 38694 23992 38700
rect 23952 38554 23980 38694
rect 23940 38548 23992 38554
rect 23940 38490 23992 38496
rect 24412 38486 24440 38830
rect 24400 38480 24452 38486
rect 24400 38422 24452 38428
rect 24584 38412 24636 38418
rect 24584 38354 24636 38360
rect 24492 38344 24544 38350
rect 24492 38286 24544 38292
rect 24504 37874 24532 38286
rect 24596 38010 24624 38354
rect 24688 38010 24716 38830
rect 24584 38004 24636 38010
rect 24584 37946 24636 37952
rect 24676 38004 24728 38010
rect 24676 37946 24728 37952
rect 24492 37868 24544 37874
rect 24492 37810 24544 37816
rect 23388 37460 23440 37466
rect 23388 37402 23440 37408
rect 24504 36922 24532 37810
rect 24492 36916 24544 36922
rect 24492 36858 24544 36864
rect 23204 36644 23256 36650
rect 23204 36586 23256 36592
rect 24964 36394 24992 41006
rect 25056 39438 25084 41414
rect 25412 40520 25464 40526
rect 25412 40462 25464 40468
rect 25424 40186 25452 40462
rect 25504 40452 25556 40458
rect 25504 40394 25556 40400
rect 25516 40186 25544 40394
rect 25412 40180 25464 40186
rect 25412 40122 25464 40128
rect 25504 40180 25556 40186
rect 25504 40122 25556 40128
rect 25424 39982 25452 40122
rect 25412 39976 25464 39982
rect 25412 39918 25464 39924
rect 25516 39438 25544 40122
rect 25044 39432 25096 39438
rect 25044 39374 25096 39380
rect 25504 39432 25556 39438
rect 25504 39374 25556 39380
rect 25044 38344 25096 38350
rect 25044 38286 25096 38292
rect 25056 37874 25084 38286
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25044 37868 25096 37874
rect 25044 37810 25096 37816
rect 25516 37670 25544 38150
rect 25504 37664 25556 37670
rect 25504 37606 25556 37612
rect 25136 36576 25188 36582
rect 25136 36518 25188 36524
rect 26068 36530 26096 43250
rect 26252 42226 26280 43318
rect 26332 43308 26384 43314
rect 26332 43250 26384 43256
rect 26344 42226 26372 43250
rect 26240 42220 26292 42226
rect 26240 42162 26292 42168
rect 26332 42220 26384 42226
rect 26332 42162 26384 42168
rect 26436 41070 26464 46378
rect 26988 45898 27016 46854
rect 27172 46510 27200 46990
rect 27620 46980 27672 46986
rect 27620 46922 27672 46928
rect 27632 46714 27660 46922
rect 27620 46708 27672 46714
rect 27620 46650 27672 46656
rect 27724 46646 27752 47620
rect 27712 46640 27764 46646
rect 27712 46582 27764 46588
rect 27160 46504 27212 46510
rect 27160 46446 27212 46452
rect 27620 45960 27672 45966
rect 27620 45902 27672 45908
rect 26976 45892 27028 45898
rect 26976 45834 27028 45840
rect 26424 41064 26476 41070
rect 26424 41006 26476 41012
rect 26240 40384 26292 40390
rect 26240 40326 26292 40332
rect 26252 40050 26280 40326
rect 26240 40044 26292 40050
rect 26240 39986 26292 39992
rect 26700 38480 26752 38486
rect 26700 38422 26752 38428
rect 26516 38276 26568 38282
rect 26516 38218 26568 38224
rect 26240 37732 26292 37738
rect 26240 37674 26292 37680
rect 26148 37664 26200 37670
rect 26148 37606 26200 37612
rect 26160 37194 26188 37606
rect 26148 37188 26200 37194
rect 26148 37130 26200 37136
rect 26252 37126 26280 37674
rect 26528 37466 26556 38218
rect 26516 37460 26568 37466
rect 26516 37402 26568 37408
rect 26712 37262 26740 38422
rect 26988 38010 27016 45834
rect 27632 44470 27660 45902
rect 27712 45892 27764 45898
rect 27712 45834 27764 45840
rect 27724 45082 27752 45834
rect 27712 45076 27764 45082
rect 27712 45018 27764 45024
rect 27620 44464 27672 44470
rect 27620 44406 27672 44412
rect 28092 44010 28120 48146
rect 28264 47660 28316 47666
rect 28264 47602 28316 47608
rect 28276 46578 28304 47602
rect 28264 46572 28316 46578
rect 28264 46514 28316 46520
rect 28276 45966 28304 46514
rect 28264 45960 28316 45966
rect 28264 45902 28316 45908
rect 28276 45490 28304 45902
rect 28448 45552 28500 45558
rect 28448 45494 28500 45500
rect 28264 45484 28316 45490
rect 28264 45426 28316 45432
rect 28276 44878 28304 45426
rect 28264 44872 28316 44878
rect 28264 44814 28316 44820
rect 28000 43982 28120 44010
rect 27436 42628 27488 42634
rect 27436 42570 27488 42576
rect 27448 42226 27476 42570
rect 27436 42220 27488 42226
rect 27436 42162 27488 42168
rect 27528 42220 27580 42226
rect 27528 42162 27580 42168
rect 27540 41818 27568 42162
rect 27712 42016 27764 42022
rect 27712 41958 27764 41964
rect 27528 41812 27580 41818
rect 27528 41754 27580 41760
rect 27540 41274 27568 41754
rect 27528 41268 27580 41274
rect 27528 41210 27580 41216
rect 27620 41064 27672 41070
rect 27620 41006 27672 41012
rect 27632 40050 27660 41006
rect 27620 40044 27672 40050
rect 27620 39986 27672 39992
rect 27528 39840 27580 39846
rect 27528 39782 27580 39788
rect 27540 39438 27568 39782
rect 27528 39432 27580 39438
rect 27528 39374 27580 39380
rect 27540 38486 27568 39374
rect 27632 39302 27660 39986
rect 27620 39296 27672 39302
rect 27620 39238 27672 39244
rect 27632 38962 27660 39238
rect 27620 38956 27672 38962
rect 27620 38898 27672 38904
rect 27724 38486 27752 41958
rect 28000 41682 28028 43982
rect 28080 42696 28132 42702
rect 28080 42638 28132 42644
rect 28092 41818 28120 42638
rect 28264 42220 28316 42226
rect 28264 42162 28316 42168
rect 28080 41812 28132 41818
rect 28080 41754 28132 41760
rect 27988 41676 28040 41682
rect 27988 41618 28040 41624
rect 28000 40594 28028 41618
rect 27988 40588 28040 40594
rect 27988 40530 28040 40536
rect 27896 40384 27948 40390
rect 27896 40326 27948 40332
rect 27908 39438 27936 40326
rect 27896 39432 27948 39438
rect 27896 39374 27948 39380
rect 27528 38480 27580 38486
rect 27528 38422 27580 38428
rect 27712 38480 27764 38486
rect 27712 38422 27764 38428
rect 26976 38004 27028 38010
rect 26976 37946 27028 37952
rect 28172 38004 28224 38010
rect 28172 37946 28224 37952
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 26700 37256 26752 37262
rect 26700 37198 26752 37204
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 26332 36712 26384 36718
rect 26332 36654 26384 36660
rect 24872 36366 24992 36394
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 24124 33856 24176 33862
rect 24124 33798 24176 33804
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 24136 33522 24164 33798
rect 24872 33522 24900 36366
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 25056 35698 25084 36110
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 25056 35290 25084 35634
rect 25044 35284 25096 35290
rect 25044 35226 25096 35232
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24032 33448 24084 33454
rect 24032 33390 24084 33396
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23860 32910 23888 33254
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 24044 32434 24072 33390
rect 24952 33380 25004 33386
rect 24952 33322 25004 33328
rect 24964 32502 24992 33322
rect 25056 32910 25084 35226
rect 25148 35086 25176 36518
rect 26068 36502 26188 36530
rect 26056 36100 26108 36106
rect 26056 36042 26108 36048
rect 25504 36032 25556 36038
rect 25504 35974 25556 35980
rect 25516 35680 25544 35974
rect 26068 35834 26096 36042
rect 26056 35828 26108 35834
rect 26056 35770 26108 35776
rect 25596 35692 25648 35698
rect 25516 35652 25596 35680
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 25516 34066 25544 35652
rect 25596 35634 25648 35640
rect 25504 34060 25556 34066
rect 25504 34002 25556 34008
rect 26056 33924 26108 33930
rect 26056 33866 26108 33872
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 25056 32570 25084 32846
rect 26068 32774 26096 33866
rect 26056 32768 26108 32774
rect 26056 32710 26108 32716
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 24952 32496 25004 32502
rect 24952 32438 25004 32444
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 25056 31890 25084 32506
rect 25136 32428 25188 32434
rect 25136 32370 25188 32376
rect 25044 31884 25096 31890
rect 25044 31826 25096 31832
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 25148 31482 25176 32370
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25504 32224 25556 32230
rect 25504 32166 25556 32172
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 25240 31346 25268 32166
rect 25516 31754 25544 32166
rect 25504 31748 25556 31754
rect 25504 31690 25556 31696
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24596 29646 24624 30194
rect 26068 30054 26096 32710
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 24596 29170 24624 29582
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 25228 29096 25280 29102
rect 25228 29038 25280 29044
rect 25240 28762 25268 29038
rect 25228 28756 25280 28762
rect 25228 28698 25280 28704
rect 26160 28558 26188 36502
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26252 35766 26280 35974
rect 26240 35760 26292 35766
rect 26240 35702 26292 35708
rect 26344 35222 26372 36654
rect 26608 36576 26660 36582
rect 26608 36518 26660 36524
rect 26620 36378 26648 36518
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26620 35562 26648 36314
rect 26700 36168 26752 36174
rect 26700 36110 26752 36116
rect 26608 35556 26660 35562
rect 26608 35498 26660 35504
rect 26712 35494 26740 36110
rect 26700 35488 26752 35494
rect 26700 35430 26752 35436
rect 26332 35216 26384 35222
rect 26332 35158 26384 35164
rect 26344 33658 26372 35158
rect 26332 33652 26384 33658
rect 26332 33594 26384 33600
rect 26240 33516 26292 33522
rect 26240 33458 26292 33464
rect 26252 32570 26280 33458
rect 26332 33380 26384 33386
rect 26332 33322 26384 33328
rect 26344 33114 26372 33322
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 26712 32978 26740 35430
rect 27264 35086 27292 37402
rect 27804 36576 27856 36582
rect 27804 36518 27856 36524
rect 27816 36174 27844 36518
rect 27528 36168 27580 36174
rect 27528 36110 27580 36116
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 27540 35290 27568 36110
rect 27528 35284 27580 35290
rect 27528 35226 27580 35232
rect 28184 35154 28212 37946
rect 28172 35148 28224 35154
rect 28172 35090 28224 35096
rect 27252 35080 27304 35086
rect 27252 35022 27304 35028
rect 27620 35080 27672 35086
rect 27620 35022 27672 35028
rect 27632 34542 27660 35022
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 27620 34536 27672 34542
rect 27620 34478 27672 34484
rect 26884 33924 26936 33930
rect 26884 33866 26936 33872
rect 26896 33454 26924 33866
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27540 33590 27568 33798
rect 27528 33584 27580 33590
rect 27528 33526 27580 33532
rect 26884 33448 26936 33454
rect 26884 33390 26936 33396
rect 26976 33448 27028 33454
rect 26976 33390 27028 33396
rect 26896 32978 26924 33390
rect 26988 32978 27016 33390
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 26700 32972 26752 32978
rect 26700 32914 26752 32920
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 26976 32972 27028 32978
rect 26976 32914 27028 32920
rect 26240 32564 26292 32570
rect 26240 32506 26292 32512
rect 26252 31414 26280 32506
rect 26988 31822 27016 32914
rect 27172 32434 27200 33254
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 27632 32366 27660 34478
rect 27712 34400 27764 34406
rect 27712 34342 27764 34348
rect 27724 33998 27752 34342
rect 28184 34202 28212 34546
rect 28172 34196 28224 34202
rect 28172 34138 28224 34144
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27988 32768 28040 32774
rect 27988 32710 28040 32716
rect 27620 32360 27672 32366
rect 27620 32302 27672 32308
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26240 31408 26292 31414
rect 26240 31350 26292 31356
rect 26988 30258 27016 31758
rect 27632 31346 27660 32302
rect 28000 31958 28028 32710
rect 27988 31952 28040 31958
rect 27988 31894 28040 31900
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27712 31136 27764 31142
rect 27712 31078 27764 31084
rect 27724 30734 27752 31078
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 27528 30592 27580 30598
rect 27528 30534 27580 30540
rect 27540 30326 27568 30534
rect 27528 30320 27580 30326
rect 27528 30262 27580 30268
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 26988 29170 27016 30194
rect 28000 29714 28028 31894
rect 28172 31340 28224 31346
rect 28172 31282 28224 31288
rect 28184 30938 28212 31282
rect 28172 30932 28224 30938
rect 28172 30874 28224 30880
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 28092 29714 28120 30194
rect 27988 29708 28040 29714
rect 27988 29650 28040 29656
rect 28080 29708 28132 29714
rect 28080 29650 28132 29656
rect 27344 29572 27396 29578
rect 27344 29514 27396 29520
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 27252 29164 27304 29170
rect 27252 29106 27304 29112
rect 27264 28762 27292 29106
rect 27252 28756 27304 28762
rect 27252 28698 27304 28704
rect 27356 28558 27384 29514
rect 28092 29306 28120 29650
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 28276 28762 28304 42162
rect 28356 40928 28408 40934
rect 28356 40870 28408 40876
rect 28368 40526 28396 40870
rect 28356 40520 28408 40526
rect 28356 40462 28408 40468
rect 28356 30592 28408 30598
rect 28356 30534 28408 30540
rect 28368 30394 28396 30534
rect 28356 30388 28408 30394
rect 28356 30330 28408 30336
rect 28368 29646 28396 30330
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28264 28756 28316 28762
rect 28264 28698 28316 28704
rect 26148 28552 26200 28558
rect 26148 28494 26200 28500
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 24872 26382 24900 28358
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 12452 19378 12480 19722
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 17420 17202 17448 21490
rect 19444 20942 19472 21490
rect 20272 21486 20300 26318
rect 26976 25832 27028 25838
rect 26976 25774 27028 25780
rect 20260 21480 20312 21486
rect 20260 21422 20312 21428
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 19854 19380 20742
rect 19444 20466 19472 20878
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19444 19854 19472 20402
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19444 19378 19472 19790
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 20088 17202 20116 19314
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 3602 9628 4422
rect 14844 4146 14872 12174
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 15304 3602 15332 3878
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9048 2650 9076 2926
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9692 800 9720 3538
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 2650 9812 3402
rect 12268 3126 12296 3470
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12544 3058 12572 3470
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 3126 12756 3334
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 15120 3058 15148 3470
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 12912 800 12940 2926
rect 15488 800 15516 3402
rect 16684 3058 16712 3878
rect 17420 3534 17448 17138
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 20272 7410 20300 21422
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 20364 10198 20392 20334
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20456 6798 20484 19722
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22480 3738 22508 4082
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16868 3126 16896 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 20364 3058 20392 3470
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16132 800 16160 2926
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 20640 800 20668 3538
rect 22848 3534 22876 4558
rect 26988 4146 27016 25774
rect 27172 9926 27200 28494
rect 28460 20942 28488 45494
rect 28552 41682 28580 51046
rect 28828 50930 28856 51206
rect 29012 51082 29040 51954
rect 28920 51054 29040 51082
rect 29196 51074 29224 54198
rect 29564 53582 29592 54606
rect 29644 54596 29696 54602
rect 29644 54538 29696 54544
rect 29656 54330 29684 54538
rect 29644 54324 29696 54330
rect 29644 54266 29696 54272
rect 29644 53984 29696 53990
rect 29644 53926 29696 53932
rect 29656 53582 29684 53926
rect 29552 53576 29604 53582
rect 29552 53518 29604 53524
rect 29644 53576 29696 53582
rect 29644 53518 29696 53524
rect 29564 52018 29592 53518
rect 30196 52488 30248 52494
rect 30196 52430 30248 52436
rect 29552 52012 29604 52018
rect 29552 51954 29604 51960
rect 29644 51400 29696 51406
rect 29644 51342 29696 51348
rect 29736 51400 29788 51406
rect 29736 51342 29788 51348
rect 28920 50998 28948 51054
rect 29196 51046 29316 51074
rect 28908 50992 28960 50998
rect 28908 50934 28960 50940
rect 28816 50924 28868 50930
rect 28816 50866 28868 50872
rect 29288 49842 29316 51046
rect 29460 50992 29512 50998
rect 29460 50934 29512 50940
rect 29092 49836 29144 49842
rect 29092 49778 29144 49784
rect 29276 49836 29328 49842
rect 29276 49778 29328 49784
rect 29000 48612 29052 48618
rect 29000 48554 29052 48560
rect 28908 47592 28960 47598
rect 28908 47534 28960 47540
rect 28816 44804 28868 44810
rect 28816 44746 28868 44752
rect 28540 41676 28592 41682
rect 28540 41618 28592 41624
rect 28552 38350 28580 41618
rect 28540 38344 28592 38350
rect 28540 38286 28592 38292
rect 28632 36712 28684 36718
rect 28632 36654 28684 36660
rect 28644 36038 28672 36654
rect 28632 36032 28684 36038
rect 28632 35974 28684 35980
rect 28644 34066 28672 35974
rect 28632 34060 28684 34066
rect 28632 34002 28684 34008
rect 28540 32836 28592 32842
rect 28540 32778 28592 32784
rect 28552 32026 28580 32778
rect 28724 32224 28776 32230
rect 28724 32166 28776 32172
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28736 31822 28764 32166
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28828 31754 28856 44746
rect 28920 43353 28948 47534
rect 29012 46170 29040 48554
rect 29000 46164 29052 46170
rect 29000 46106 29052 46112
rect 29000 45416 29052 45422
rect 29000 45358 29052 45364
rect 29012 45014 29040 45358
rect 29000 45008 29052 45014
rect 29000 44950 29052 44956
rect 29104 44878 29132 49778
rect 29184 49428 29236 49434
rect 29184 49370 29236 49376
rect 29196 48618 29224 49370
rect 29184 48612 29236 48618
rect 29184 48554 29236 48560
rect 29288 48142 29316 49778
rect 29472 49434 29500 50934
rect 29552 49972 29604 49978
rect 29552 49914 29604 49920
rect 29460 49428 29512 49434
rect 29460 49370 29512 49376
rect 29564 49230 29592 49914
rect 29552 49224 29604 49230
rect 29552 49166 29604 49172
rect 29368 48816 29420 48822
rect 29420 48764 29500 48770
rect 29368 48760 29500 48764
rect 29368 48758 29512 48760
rect 29380 48754 29512 48758
rect 29380 48742 29460 48754
rect 29460 48696 29512 48702
rect 29564 48618 29592 49166
rect 29656 48822 29684 51342
rect 29748 50726 29776 51342
rect 29828 50788 29880 50794
rect 29828 50730 29880 50736
rect 29736 50720 29788 50726
rect 29736 50662 29788 50668
rect 29748 49298 29776 50662
rect 29840 50318 29868 50730
rect 29828 50312 29880 50318
rect 29828 50254 29880 50260
rect 30012 50312 30064 50318
rect 30012 50254 30064 50260
rect 30208 50300 30236 52430
rect 30472 52012 30524 52018
rect 30472 51954 30524 51960
rect 31392 52012 31444 52018
rect 31392 51954 31444 51960
rect 30484 51610 30512 51954
rect 30472 51604 30524 51610
rect 30472 51546 30524 51552
rect 31404 51406 31432 51954
rect 31392 51400 31444 51406
rect 31392 51342 31444 51348
rect 31404 50930 31432 51342
rect 31392 50924 31444 50930
rect 31392 50866 31444 50872
rect 30840 50720 30892 50726
rect 30840 50662 30892 50668
rect 30852 50386 30880 50662
rect 30840 50380 30892 50386
rect 30840 50322 30892 50328
rect 30288 50312 30340 50318
rect 30208 50272 30288 50300
rect 29920 50176 29972 50182
rect 29920 50118 29972 50124
rect 29932 49434 29960 50118
rect 29920 49428 29972 49434
rect 29920 49370 29972 49376
rect 29736 49292 29788 49298
rect 29736 49234 29788 49240
rect 29644 48816 29696 48822
rect 29644 48758 29696 48764
rect 29552 48612 29604 48618
rect 29552 48554 29604 48560
rect 29276 48136 29328 48142
rect 29276 48078 29328 48084
rect 29552 47728 29604 47734
rect 29552 47670 29604 47676
rect 29276 45008 29328 45014
rect 29276 44950 29328 44956
rect 29092 44872 29144 44878
rect 29092 44814 29144 44820
rect 29104 43858 29132 44814
rect 29092 43852 29144 43858
rect 29092 43794 29144 43800
rect 29092 43716 29144 43722
rect 29092 43658 29144 43664
rect 28906 43344 28962 43353
rect 28906 43279 28962 43288
rect 29000 42696 29052 42702
rect 29000 42638 29052 42644
rect 29012 41818 29040 42638
rect 29000 41812 29052 41818
rect 29000 41754 29052 41760
rect 28908 41608 28960 41614
rect 28908 41550 28960 41556
rect 29000 41608 29052 41614
rect 29000 41550 29052 41556
rect 28920 39914 28948 41550
rect 28908 39908 28960 39914
rect 28908 39850 28960 39856
rect 29012 39846 29040 41550
rect 29000 39840 29052 39846
rect 29000 39782 29052 39788
rect 28908 39500 28960 39506
rect 28908 39442 28960 39448
rect 28920 39098 28948 39442
rect 29104 39098 29132 43658
rect 29288 41414 29316 44950
rect 29460 44396 29512 44402
rect 29460 44338 29512 44344
rect 29472 43994 29500 44338
rect 29460 43988 29512 43994
rect 29460 43930 29512 43936
rect 29368 42560 29420 42566
rect 29368 42502 29420 42508
rect 29460 42560 29512 42566
rect 29460 42502 29512 42508
rect 29380 41682 29408 42502
rect 29472 41970 29500 42502
rect 29564 42362 29592 47670
rect 30024 47190 30052 50254
rect 30104 50244 30156 50250
rect 30104 50186 30156 50192
rect 30116 49978 30144 50186
rect 30104 49972 30156 49978
rect 30104 49914 30156 49920
rect 30104 49768 30156 49774
rect 30104 49710 30156 49716
rect 30116 49230 30144 49710
rect 30104 49224 30156 49230
rect 30104 49166 30156 49172
rect 30208 48278 30236 50272
rect 30288 50254 30340 50260
rect 30932 50312 30984 50318
rect 30932 50254 30984 50260
rect 30944 49978 30972 50254
rect 30932 49972 30984 49978
rect 30932 49914 30984 49920
rect 30564 49156 30616 49162
rect 30564 49098 30616 49104
rect 30196 48272 30248 48278
rect 30196 48214 30248 48220
rect 30472 48068 30524 48074
rect 30472 48010 30524 48016
rect 30380 47660 30432 47666
rect 30380 47602 30432 47608
rect 30012 47184 30064 47190
rect 30012 47126 30064 47132
rect 30288 47184 30340 47190
rect 30288 47126 30340 47132
rect 30104 47116 30156 47122
rect 30104 47058 30156 47064
rect 30012 46708 30064 46714
rect 30012 46650 30064 46656
rect 29920 46504 29972 46510
rect 29920 46446 29972 46452
rect 29932 46374 29960 46446
rect 29920 46368 29972 46374
rect 29920 46310 29972 46316
rect 29736 46028 29788 46034
rect 29736 45970 29788 45976
rect 29552 42356 29604 42362
rect 29552 42298 29604 42304
rect 29564 42242 29592 42298
rect 29564 42214 29684 42242
rect 29472 41942 29592 41970
rect 29368 41676 29420 41682
rect 29368 41618 29420 41624
rect 29288 41386 29500 41414
rect 29276 41200 29328 41206
rect 29276 41142 29328 41148
rect 29184 40996 29236 41002
rect 29184 40938 29236 40944
rect 28908 39092 28960 39098
rect 28908 39034 28960 39040
rect 29092 39092 29144 39098
rect 29092 39034 29144 39040
rect 29000 36712 29052 36718
rect 29196 36666 29224 40938
rect 29288 38434 29316 41142
rect 29368 40112 29420 40118
rect 29368 40054 29420 40060
rect 29380 38554 29408 40054
rect 29368 38548 29420 38554
rect 29368 38490 29420 38496
rect 29288 38406 29408 38434
rect 29380 36786 29408 38406
rect 29368 36780 29420 36786
rect 29368 36722 29420 36728
rect 29000 36654 29052 36660
rect 29012 35698 29040 36654
rect 29104 36638 29224 36666
rect 29276 36712 29328 36718
rect 29276 36654 29328 36660
rect 29000 35692 29052 35698
rect 29000 35634 29052 35640
rect 29104 35578 29132 36638
rect 29104 35550 29224 35578
rect 29092 33856 29144 33862
rect 29092 33798 29144 33804
rect 29104 33318 29132 33798
rect 29092 33312 29144 33318
rect 29092 33254 29144 33260
rect 29000 32768 29052 32774
rect 29000 32710 29052 32716
rect 28828 31726 28948 31754
rect 28816 31272 28868 31278
rect 28816 31214 28868 31220
rect 28828 30258 28856 31214
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 28540 29504 28592 29510
rect 28540 29446 28592 29452
rect 28552 28626 28580 29446
rect 28540 28620 28592 28626
rect 28540 28562 28592 28568
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28828 27674 28856 28018
rect 28816 27668 28868 27674
rect 28816 27610 28868 27616
rect 28724 27396 28776 27402
rect 28724 27338 28776 27344
rect 28736 26976 28764 27338
rect 28736 26948 28856 26976
rect 28828 26858 28856 26948
rect 28816 26852 28868 26858
rect 28816 26794 28868 26800
rect 28828 26314 28856 26794
rect 28816 26308 28868 26314
rect 28816 26250 28868 26256
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 28920 6914 28948 31726
rect 29012 31482 29040 32710
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 29012 28558 29040 31078
rect 29104 30054 29132 33254
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 29012 28014 29040 28494
rect 29000 28008 29052 28014
rect 29052 27956 29132 27962
rect 29000 27950 29132 27956
rect 29012 27934 29132 27950
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 29012 26926 29040 27814
rect 29104 27470 29132 27934
rect 29092 27464 29144 27470
rect 29092 27406 29144 27412
rect 29000 26920 29052 26926
rect 29000 26862 29052 26868
rect 28828 6886 28948 6914
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 23032 3126 23060 3878
rect 23308 3194 23336 3878
rect 26896 3602 26924 3878
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23204 2984 23256 2990
rect 23204 2926 23256 2932
rect 23216 800 23244 2926
rect 25148 800 25176 3538
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26712 3058 26740 3470
rect 26988 3398 27016 4082
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 26976 3392 27028 3398
rect 26976 3334 27028 3340
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 27080 800 27108 3538
rect 28828 3466 28856 6886
rect 29196 4078 29224 35550
rect 29288 35494 29316 36654
rect 29276 35488 29328 35494
rect 29276 35430 29328 35436
rect 29288 30734 29316 35430
rect 29276 30728 29328 30734
rect 29276 30670 29328 30676
rect 29276 28076 29328 28082
rect 29276 28018 29328 28024
rect 29288 27878 29316 28018
rect 29368 27940 29420 27946
rect 29368 27882 29420 27888
rect 29276 27872 29328 27878
rect 29276 27814 29328 27820
rect 29276 27532 29328 27538
rect 29380 27520 29408 27882
rect 29328 27492 29408 27520
rect 29276 27474 29328 27480
rect 29380 26382 29408 27492
rect 29368 26376 29420 26382
rect 29368 26318 29420 26324
rect 29368 25696 29420 25702
rect 29368 25638 29420 25644
rect 29380 10062 29408 25638
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 29472 6322 29500 41386
rect 29564 41138 29592 41942
rect 29552 41132 29604 41138
rect 29552 41074 29604 41080
rect 29552 38956 29604 38962
rect 29552 38898 29604 38904
rect 29564 38010 29592 38898
rect 29552 38004 29604 38010
rect 29552 37946 29604 37952
rect 29656 37262 29684 42214
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 29656 36854 29684 37198
rect 29644 36848 29696 36854
rect 29644 36790 29696 36796
rect 29552 32768 29604 32774
rect 29552 32710 29604 32716
rect 29564 32434 29592 32710
rect 29552 32428 29604 32434
rect 29552 32370 29604 32376
rect 29748 31754 29776 45970
rect 29932 45370 29960 46310
rect 30024 45558 30052 46650
rect 30012 45552 30064 45558
rect 30012 45494 30064 45500
rect 29932 45342 30052 45370
rect 29828 42220 29880 42226
rect 29828 42162 29880 42168
rect 29840 41138 29868 42162
rect 29920 41744 29972 41750
rect 29920 41686 29972 41692
rect 29828 41132 29880 41138
rect 29828 41074 29880 41080
rect 29840 39574 29868 41074
rect 29932 40730 29960 41686
rect 30024 41002 30052 45342
rect 30012 40996 30064 41002
rect 30012 40938 30064 40944
rect 29920 40724 29972 40730
rect 29920 40666 29972 40672
rect 30116 40594 30144 47058
rect 30300 46578 30328 47126
rect 30288 46572 30340 46578
rect 30288 46514 30340 46520
rect 30392 46034 30420 47602
rect 30484 47598 30512 48010
rect 30576 47734 30604 49098
rect 31024 48136 31076 48142
rect 31024 48078 31076 48084
rect 30564 47728 30616 47734
rect 30564 47670 30616 47676
rect 30472 47592 30524 47598
rect 30472 47534 30524 47540
rect 30484 46900 30512 47534
rect 30576 47054 30604 47670
rect 31036 47190 31064 48078
rect 31024 47184 31076 47190
rect 31024 47126 31076 47132
rect 30656 47116 30708 47122
rect 30656 47058 30708 47064
rect 30564 47048 30616 47054
rect 30564 46990 30616 46996
rect 30484 46872 30604 46900
rect 30380 46028 30432 46034
rect 30380 45970 30432 45976
rect 30288 44872 30340 44878
rect 30288 44814 30340 44820
rect 30196 44192 30248 44198
rect 30196 44134 30248 44140
rect 30208 42702 30236 44134
rect 30196 42696 30248 42702
rect 30196 42638 30248 42644
rect 30208 41138 30236 42638
rect 30196 41132 30248 41138
rect 30196 41074 30248 41080
rect 30196 40996 30248 41002
rect 30196 40938 30248 40944
rect 30104 40588 30156 40594
rect 30024 40548 30104 40576
rect 29828 39568 29880 39574
rect 29828 39510 29880 39516
rect 29840 39098 29868 39510
rect 29828 39092 29880 39098
rect 29828 39034 29880 39040
rect 29840 38214 29868 39034
rect 30024 38962 30052 40548
rect 30104 40530 30156 40536
rect 30208 40186 30236 40938
rect 30196 40180 30248 40186
rect 30196 40122 30248 40128
rect 30208 39438 30236 40122
rect 30300 39914 30328 44814
rect 30472 42152 30524 42158
rect 30472 42094 30524 42100
rect 30380 42016 30432 42022
rect 30380 41958 30432 41964
rect 30392 40390 30420 41958
rect 30484 41138 30512 42094
rect 30472 41132 30524 41138
rect 30472 41074 30524 41080
rect 30484 40390 30512 41074
rect 30380 40384 30432 40390
rect 30380 40326 30432 40332
rect 30472 40384 30524 40390
rect 30472 40326 30524 40332
rect 30392 40186 30420 40326
rect 30380 40180 30432 40186
rect 30380 40122 30432 40128
rect 30392 40050 30420 40122
rect 30380 40044 30432 40050
rect 30380 39986 30432 39992
rect 30288 39908 30340 39914
rect 30288 39850 30340 39856
rect 30196 39432 30248 39438
rect 30196 39374 30248 39380
rect 30288 39296 30340 39302
rect 30288 39238 30340 39244
rect 30012 38956 30064 38962
rect 30012 38898 30064 38904
rect 30196 38956 30248 38962
rect 30196 38898 30248 38904
rect 30024 38758 30052 38898
rect 30012 38752 30064 38758
rect 30012 38694 30064 38700
rect 29828 38208 29880 38214
rect 29828 38150 29880 38156
rect 30024 37806 30052 38694
rect 30104 38276 30156 38282
rect 30104 38218 30156 38224
rect 30116 37806 30144 38218
rect 30208 37942 30236 38898
rect 30300 38486 30328 39238
rect 30484 39030 30512 40326
rect 30472 39024 30524 39030
rect 30472 38966 30524 38972
rect 30288 38480 30340 38486
rect 30288 38422 30340 38428
rect 30196 37936 30248 37942
rect 30196 37878 30248 37884
rect 30012 37800 30064 37806
rect 30012 37742 30064 37748
rect 30104 37800 30156 37806
rect 30104 37742 30156 37748
rect 30024 37262 30052 37742
rect 30012 37256 30064 37262
rect 30012 37198 30064 37204
rect 30300 37194 30328 38422
rect 30484 38350 30512 38966
rect 30380 38344 30432 38350
rect 30380 38286 30432 38292
rect 30472 38344 30524 38350
rect 30472 38286 30524 38292
rect 30392 37466 30420 38286
rect 30484 38010 30512 38286
rect 30472 38004 30524 38010
rect 30472 37946 30524 37952
rect 30380 37460 30432 37466
rect 30380 37402 30432 37408
rect 30288 37188 30340 37194
rect 30288 37130 30340 37136
rect 29828 36576 29880 36582
rect 29828 36518 29880 36524
rect 30472 36576 30524 36582
rect 30472 36518 30524 36524
rect 29840 36242 29868 36518
rect 29828 36236 29880 36242
rect 29828 36178 29880 36184
rect 30380 35760 30432 35766
rect 30380 35702 30432 35708
rect 30012 35284 30064 35290
rect 30012 35226 30064 35232
rect 29920 33856 29972 33862
rect 29920 33798 29972 33804
rect 29932 33590 29960 33798
rect 29920 33584 29972 33590
rect 29920 33526 29972 33532
rect 29932 33046 29960 33526
rect 29920 33040 29972 33046
rect 29920 32982 29972 32988
rect 30024 32978 30052 35226
rect 30104 34944 30156 34950
rect 30104 34886 30156 34892
rect 30116 34066 30144 34886
rect 30392 34678 30420 35702
rect 30380 34672 30432 34678
rect 30380 34614 30432 34620
rect 30392 34066 30420 34614
rect 30104 34060 30156 34066
rect 30104 34002 30156 34008
rect 30380 34060 30432 34066
rect 30380 34002 30432 34008
rect 30116 33590 30144 34002
rect 30104 33584 30156 33590
rect 30104 33526 30156 33532
rect 30012 32972 30064 32978
rect 30012 32914 30064 32920
rect 30288 32972 30340 32978
rect 30288 32914 30340 32920
rect 29748 31726 29960 31754
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 29550 27568 29606 27577
rect 29550 27503 29606 27512
rect 29564 26994 29592 27503
rect 29552 26988 29604 26994
rect 29552 26930 29604 26936
rect 29564 25838 29592 26930
rect 29656 26926 29684 27950
rect 29840 27946 29868 28494
rect 29828 27940 29880 27946
rect 29828 27882 29880 27888
rect 29828 27396 29880 27402
rect 29828 27338 29880 27344
rect 29840 27130 29868 27338
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 29644 26920 29696 26926
rect 29644 26862 29696 26868
rect 29748 26382 29776 26930
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29552 25832 29604 25838
rect 29552 25774 29604 25780
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29656 20874 29684 21490
rect 29644 20868 29696 20874
rect 29644 20810 29696 20816
rect 29656 20466 29684 20810
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29656 19854 29684 20402
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29656 19378 29684 19790
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29552 16652 29604 16658
rect 29552 16594 29604 16600
rect 29564 9586 29592 16594
rect 29736 9988 29788 9994
rect 29736 9930 29788 9936
rect 29748 9722 29776 9930
rect 29736 9716 29788 9722
rect 29736 9658 29788 9664
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29932 6914 29960 31726
rect 30300 31278 30328 32914
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30392 31890 30420 32302
rect 30380 31884 30432 31890
rect 30380 31826 30432 31832
rect 30484 31754 30512 36518
rect 30392 31726 30512 31754
rect 30288 31272 30340 31278
rect 30288 31214 30340 31220
rect 30196 31136 30248 31142
rect 30196 31078 30248 31084
rect 30208 30666 30236 31078
rect 30300 30802 30328 31214
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30196 30660 30248 30666
rect 30196 30602 30248 30608
rect 30392 28490 30420 31726
rect 30472 30048 30524 30054
rect 30472 29990 30524 29996
rect 30484 29578 30512 29990
rect 30472 29572 30524 29578
rect 30472 29514 30524 29520
rect 30484 29170 30512 29514
rect 30472 29164 30524 29170
rect 30472 29106 30524 29112
rect 30380 28484 30432 28490
rect 30380 28426 30432 28432
rect 30472 27464 30524 27470
rect 30472 27406 30524 27412
rect 30288 27396 30340 27402
rect 30288 27338 30340 27344
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 30024 26382 30052 26862
rect 30300 26382 30328 27338
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30012 26376 30064 26382
rect 30288 26376 30340 26382
rect 30012 26318 30064 26324
rect 30194 26344 30250 26353
rect 30288 26318 30340 26324
rect 30194 26279 30196 26288
rect 30248 26279 30250 26288
rect 30196 26250 30248 26256
rect 30392 25906 30420 27270
rect 30484 27062 30512 27406
rect 30472 27056 30524 27062
rect 30472 26998 30524 27004
rect 30380 25900 30432 25906
rect 30380 25842 30432 25848
rect 30576 22094 30604 46872
rect 30668 36582 30696 47058
rect 31036 46646 31064 47126
rect 31392 46980 31444 46986
rect 31392 46922 31444 46928
rect 31404 46714 31432 46922
rect 31392 46708 31444 46714
rect 31392 46650 31444 46656
rect 31024 46640 31076 46646
rect 31024 46582 31076 46588
rect 31036 46034 31064 46582
rect 31024 46028 31076 46034
rect 31024 45970 31076 45976
rect 31036 45422 31064 45970
rect 31024 45416 31076 45422
rect 31024 45358 31076 45364
rect 31036 45082 31064 45358
rect 31024 45076 31076 45082
rect 31024 45018 31076 45024
rect 31036 44470 31064 45018
rect 31024 44464 31076 44470
rect 31024 44406 31076 44412
rect 31036 43858 31064 44406
rect 31024 43852 31076 43858
rect 31024 43794 31076 43800
rect 30932 42764 30984 42770
rect 30932 42706 30984 42712
rect 30840 41268 30892 41274
rect 30840 41210 30892 41216
rect 30748 40928 30800 40934
rect 30748 40870 30800 40876
rect 30760 39098 30788 40870
rect 30852 40050 30880 41210
rect 30840 40044 30892 40050
rect 30840 39986 30892 39992
rect 30748 39092 30800 39098
rect 30748 39034 30800 39040
rect 30840 38956 30892 38962
rect 30944 38944 30972 42706
rect 31300 42696 31352 42702
rect 31300 42638 31352 42644
rect 31208 42016 31260 42022
rect 31208 41958 31260 41964
rect 31220 41857 31248 41958
rect 31206 41848 31262 41857
rect 31312 41818 31340 42638
rect 31392 42220 31444 42226
rect 31392 42162 31444 42168
rect 31206 41783 31262 41792
rect 31300 41812 31352 41818
rect 31300 41754 31352 41760
rect 31208 41744 31260 41750
rect 31208 41686 31260 41692
rect 31116 41540 31168 41546
rect 31116 41482 31168 41488
rect 31128 40458 31156 41482
rect 31116 40452 31168 40458
rect 31116 40394 31168 40400
rect 31024 39092 31076 39098
rect 31024 39034 31076 39040
rect 30892 38916 30972 38944
rect 30840 38898 30892 38904
rect 30748 38344 30800 38350
rect 30748 38286 30800 38292
rect 30760 37874 30788 38286
rect 30748 37868 30800 37874
rect 30748 37810 30800 37816
rect 30656 36576 30708 36582
rect 30656 36518 30708 36524
rect 30748 35760 30800 35766
rect 30748 35702 30800 35708
rect 30760 35154 30788 35702
rect 30748 35148 30800 35154
rect 30748 35090 30800 35096
rect 30852 35086 30880 38898
rect 30932 38752 30984 38758
rect 30932 38694 30984 38700
rect 30944 38418 30972 38694
rect 30932 38412 30984 38418
rect 30932 38354 30984 38360
rect 30930 38312 30986 38321
rect 30930 38247 30986 38256
rect 30944 35766 30972 38247
rect 31036 37890 31064 39034
rect 31128 38729 31156 40394
rect 31114 38720 31170 38729
rect 31114 38655 31170 38664
rect 31116 38412 31168 38418
rect 31116 38354 31168 38360
rect 31128 38010 31156 38354
rect 31116 38004 31168 38010
rect 31116 37946 31168 37952
rect 31036 37862 31156 37890
rect 31024 37800 31076 37806
rect 31024 37742 31076 37748
rect 31036 37262 31064 37742
rect 31128 37466 31156 37862
rect 31116 37460 31168 37466
rect 31116 37402 31168 37408
rect 31220 37262 31248 41686
rect 31312 40730 31340 41754
rect 31404 41070 31432 42162
rect 31392 41064 31444 41070
rect 31392 41006 31444 41012
rect 31300 40724 31352 40730
rect 31300 40666 31352 40672
rect 31312 40118 31340 40666
rect 31404 40662 31432 41006
rect 31392 40656 31444 40662
rect 31392 40598 31444 40604
rect 31300 40112 31352 40118
rect 31300 40054 31352 40060
rect 31496 39522 31524 56374
rect 32140 56370 32168 57190
rect 32128 56364 32180 56370
rect 32128 56306 32180 56312
rect 32876 56302 32904 59200
rect 33520 57458 33548 59200
rect 33508 57452 33560 57458
rect 33508 57394 33560 57400
rect 33600 57248 33652 57254
rect 33600 57190 33652 57196
rect 35624 57248 35676 57254
rect 35624 57190 35676 57196
rect 32404 56296 32456 56302
rect 32404 56238 32456 56244
rect 32864 56296 32916 56302
rect 32864 56238 32916 56244
rect 32416 55894 32444 56238
rect 32404 55888 32456 55894
rect 32404 55830 32456 55836
rect 32220 55752 32272 55758
rect 32220 55694 32272 55700
rect 32128 52080 32180 52086
rect 32128 52022 32180 52028
rect 32140 51406 32168 52022
rect 32128 51400 32180 51406
rect 32128 51342 32180 51348
rect 32140 50862 32168 51342
rect 31668 50856 31720 50862
rect 31668 50798 31720 50804
rect 31944 50856 31996 50862
rect 31944 50798 31996 50804
rect 32128 50856 32180 50862
rect 32128 50798 32180 50804
rect 31680 49910 31708 50798
rect 31956 50522 31984 50798
rect 31944 50516 31996 50522
rect 31944 50458 31996 50464
rect 32140 50318 32168 50798
rect 32128 50312 32180 50318
rect 32128 50254 32180 50260
rect 31668 49904 31720 49910
rect 31668 49846 31720 49852
rect 32140 49230 32168 50254
rect 32128 49224 32180 49230
rect 32128 49166 32180 49172
rect 31944 48816 31996 48822
rect 31944 48758 31996 48764
rect 31956 48074 31984 48758
rect 31944 48068 31996 48074
rect 31944 48010 31996 48016
rect 31760 48000 31812 48006
rect 31760 47942 31812 47948
rect 31576 42696 31628 42702
rect 31576 42638 31628 42644
rect 31588 41546 31616 42638
rect 31576 41540 31628 41546
rect 31576 41482 31628 41488
rect 31772 40984 31800 47942
rect 31956 47666 31984 48010
rect 31944 47660 31996 47666
rect 31944 47602 31996 47608
rect 31852 47456 31904 47462
rect 31852 47398 31904 47404
rect 31864 47122 31892 47398
rect 31852 47116 31904 47122
rect 31852 47058 31904 47064
rect 31956 42770 31984 47602
rect 32128 46368 32180 46374
rect 32128 46310 32180 46316
rect 32140 45966 32168 46310
rect 32128 45960 32180 45966
rect 32128 45902 32180 45908
rect 32036 45348 32088 45354
rect 32036 45290 32088 45296
rect 32048 44946 32076 45290
rect 32036 44940 32088 44946
rect 32036 44882 32088 44888
rect 32048 44470 32076 44882
rect 32232 44878 32260 55694
rect 33612 55622 33640 57190
rect 34934 57148 35242 57168
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57072 35242 57092
rect 35636 56846 35664 57190
rect 35624 56840 35676 56846
rect 35624 56782 35676 56788
rect 36096 56778 36124 59200
rect 35808 56772 35860 56778
rect 35808 56714 35860 56720
rect 36084 56772 36136 56778
rect 36084 56714 36136 56720
rect 35716 56160 35768 56166
rect 35716 56102 35768 56108
rect 34934 56060 35242 56080
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55984 35242 56004
rect 35728 55758 35756 56102
rect 35820 55894 35848 56714
rect 35808 55888 35860 55894
rect 35808 55830 35860 55836
rect 35348 55752 35400 55758
rect 35348 55694 35400 55700
rect 35716 55752 35768 55758
rect 35716 55694 35768 55700
rect 33600 55616 33652 55622
rect 33600 55558 33652 55564
rect 34934 54972 35242 54992
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54896 35242 54916
rect 34428 54596 34480 54602
rect 34428 54538 34480 54544
rect 32404 51944 32456 51950
rect 32404 51886 32456 51892
rect 32312 51808 32364 51814
rect 32312 51750 32364 51756
rect 32324 51406 32352 51750
rect 32312 51400 32364 51406
rect 32312 51342 32364 51348
rect 32416 51218 32444 51886
rect 32588 51400 32640 51406
rect 32588 51342 32640 51348
rect 32496 51332 32548 51338
rect 32496 51274 32548 51280
rect 32324 51190 32444 51218
rect 32324 50182 32352 51190
rect 32312 50176 32364 50182
rect 32312 50118 32364 50124
rect 32324 49978 32352 50118
rect 32508 49978 32536 51274
rect 32600 51066 32628 51342
rect 33140 51332 33192 51338
rect 33140 51274 33192 51280
rect 33048 51264 33100 51270
rect 33048 51206 33100 51212
rect 32588 51060 32640 51066
rect 32588 51002 32640 51008
rect 32680 50924 32732 50930
rect 32680 50866 32732 50872
rect 32692 49978 32720 50866
rect 32312 49972 32364 49978
rect 32312 49914 32364 49920
rect 32496 49972 32548 49978
rect 32496 49914 32548 49920
rect 32680 49972 32732 49978
rect 32680 49914 32732 49920
rect 33060 49842 33088 51206
rect 33152 51066 33180 51274
rect 33416 51264 33468 51270
rect 33416 51206 33468 51212
rect 33876 51264 33928 51270
rect 33876 51206 33928 51212
rect 33428 51074 33456 51206
rect 33140 51060 33192 51066
rect 33140 51002 33192 51008
rect 33336 51046 33456 51074
rect 33336 50930 33364 51046
rect 33888 50998 33916 51206
rect 33876 50992 33928 50998
rect 33876 50934 33928 50940
rect 33324 50924 33376 50930
rect 33324 50866 33376 50872
rect 33336 50522 33364 50866
rect 33508 50856 33560 50862
rect 33508 50798 33560 50804
rect 33520 50522 33548 50798
rect 33968 50720 34020 50726
rect 33968 50662 34020 50668
rect 33324 50516 33376 50522
rect 33324 50458 33376 50464
rect 33508 50516 33560 50522
rect 33508 50458 33560 50464
rect 33140 50244 33192 50250
rect 33140 50186 33192 50192
rect 33152 49978 33180 50186
rect 33140 49972 33192 49978
rect 33140 49914 33192 49920
rect 33520 49910 33548 50458
rect 33980 50182 34008 50662
rect 33968 50176 34020 50182
rect 33968 50118 34020 50124
rect 33508 49904 33560 49910
rect 33508 49846 33560 49852
rect 33048 49836 33100 49842
rect 33048 49778 33100 49784
rect 34244 49156 34296 49162
rect 34244 49098 34296 49104
rect 34256 48890 34284 49098
rect 34244 48884 34296 48890
rect 34244 48826 34296 48832
rect 33692 48748 33744 48754
rect 33692 48690 33744 48696
rect 32588 48680 32640 48686
rect 32588 48622 32640 48628
rect 32600 47666 32628 48622
rect 33048 48068 33100 48074
rect 33048 48010 33100 48016
rect 33060 47802 33088 48010
rect 33704 48006 33732 48690
rect 34152 48136 34204 48142
rect 34152 48078 34204 48084
rect 33324 48000 33376 48006
rect 33324 47942 33376 47948
rect 33692 48000 33744 48006
rect 33692 47942 33744 47948
rect 33048 47796 33100 47802
rect 33048 47738 33100 47744
rect 33336 47666 33364 47942
rect 33876 47796 33928 47802
rect 33876 47738 33928 47744
rect 32404 47660 32456 47666
rect 32404 47602 32456 47608
rect 32588 47660 32640 47666
rect 33324 47660 33376 47666
rect 32640 47620 32720 47648
rect 32588 47602 32640 47608
rect 32416 46578 32444 47602
rect 32404 46572 32456 46578
rect 32404 46514 32456 46520
rect 32416 44878 32444 46514
rect 32588 46436 32640 46442
rect 32588 46378 32640 46384
rect 32600 45830 32628 46378
rect 32588 45824 32640 45830
rect 32588 45766 32640 45772
rect 32220 44872 32272 44878
rect 32220 44814 32272 44820
rect 32404 44872 32456 44878
rect 32404 44814 32456 44820
rect 32036 44464 32088 44470
rect 32036 44406 32088 44412
rect 32416 44402 32444 44814
rect 32404 44396 32456 44402
rect 32404 44338 32456 44344
rect 32404 44260 32456 44266
rect 32404 44202 32456 44208
rect 32128 44192 32180 44198
rect 32128 44134 32180 44140
rect 32140 43790 32168 44134
rect 32128 43784 32180 43790
rect 32128 43726 32180 43732
rect 32416 43654 32444 44202
rect 32404 43648 32456 43654
rect 32404 43590 32456 43596
rect 31944 42764 31996 42770
rect 31944 42706 31996 42712
rect 31956 42378 31984 42706
rect 32312 42560 32364 42566
rect 32312 42502 32364 42508
rect 31956 42350 32168 42378
rect 32036 42084 32088 42090
rect 32036 42026 32088 42032
rect 31944 41472 31996 41478
rect 31944 41414 31996 41420
rect 31852 40996 31904 41002
rect 31772 40956 31852 40984
rect 31772 40730 31800 40956
rect 31852 40938 31904 40944
rect 31760 40724 31812 40730
rect 31760 40666 31812 40672
rect 31772 40594 31800 40666
rect 31760 40588 31812 40594
rect 31760 40530 31812 40536
rect 31668 40520 31720 40526
rect 31668 40462 31720 40468
rect 31680 40186 31708 40462
rect 31668 40180 31720 40186
rect 31668 40122 31720 40128
rect 31852 39840 31904 39846
rect 31852 39782 31904 39788
rect 31404 39494 31524 39522
rect 31298 38720 31354 38729
rect 31298 38655 31354 38664
rect 31312 38321 31340 38655
rect 31298 38312 31354 38321
rect 31298 38247 31354 38256
rect 31300 38208 31352 38214
rect 31300 38150 31352 38156
rect 31312 37738 31340 38150
rect 31300 37732 31352 37738
rect 31300 37674 31352 37680
rect 31312 37330 31340 37674
rect 31300 37324 31352 37330
rect 31300 37266 31352 37272
rect 31024 37256 31076 37262
rect 31024 37198 31076 37204
rect 31208 37256 31260 37262
rect 31208 37198 31260 37204
rect 31036 36825 31064 37198
rect 31022 36816 31078 36825
rect 31022 36751 31078 36760
rect 31024 36168 31076 36174
rect 31024 36110 31076 36116
rect 30932 35760 30984 35766
rect 30932 35702 30984 35708
rect 30932 35216 30984 35222
rect 30932 35158 30984 35164
rect 30840 35080 30892 35086
rect 30840 35022 30892 35028
rect 30748 33924 30800 33930
rect 30748 33866 30800 33872
rect 30760 33658 30788 33866
rect 30748 33652 30800 33658
rect 30748 33594 30800 33600
rect 30944 33522 30972 35158
rect 31036 35154 31064 36110
rect 31024 35148 31076 35154
rect 31024 35090 31076 35096
rect 30932 33516 30984 33522
rect 30932 33458 30984 33464
rect 30932 31884 30984 31890
rect 30932 31826 30984 31832
rect 30944 31482 30972 31826
rect 30932 31476 30984 31482
rect 30932 31418 30984 31424
rect 31116 31340 31168 31346
rect 31116 31282 31168 31288
rect 31128 30954 31156 31282
rect 31128 30938 31248 30954
rect 31128 30932 31260 30938
rect 31128 30926 31208 30932
rect 31128 30190 31156 30926
rect 31208 30874 31260 30880
rect 31116 30184 31168 30190
rect 31116 30126 31168 30132
rect 30840 30048 30892 30054
rect 30840 29990 30892 29996
rect 30852 29782 30880 29990
rect 30840 29776 30892 29782
rect 30840 29718 30892 29724
rect 30852 29646 30880 29718
rect 31128 29714 31156 30126
rect 31116 29708 31168 29714
rect 31116 29650 31168 29656
rect 30840 29640 30892 29646
rect 30840 29582 30892 29588
rect 30852 29034 30880 29582
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 30840 29028 30892 29034
rect 30840 28970 30892 28976
rect 31036 28218 31064 29106
rect 31116 28552 31168 28558
rect 31116 28494 31168 28500
rect 31024 28212 31076 28218
rect 31024 28154 31076 28160
rect 31128 28014 31156 28494
rect 31208 28076 31260 28082
rect 31208 28018 31260 28024
rect 31116 28008 31168 28014
rect 31116 27950 31168 27956
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30760 27130 30788 27406
rect 30748 27124 30800 27130
rect 30748 27066 30800 27072
rect 31128 26994 31156 27950
rect 31116 26988 31168 26994
rect 31116 26930 31168 26936
rect 31220 26926 31248 28018
rect 31300 27532 31352 27538
rect 31300 27474 31352 27480
rect 31312 27062 31340 27474
rect 31300 27056 31352 27062
rect 31300 26998 31352 27004
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 31208 26920 31260 26926
rect 31208 26862 31260 26868
rect 31300 26920 31352 26926
rect 31300 26862 31352 26868
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30668 25906 30696 26726
rect 30852 26450 30880 26794
rect 30840 26444 30892 26450
rect 30840 26386 30892 26392
rect 30944 26382 30972 26862
rect 30748 26376 30800 26382
rect 30746 26344 30748 26353
rect 30932 26376 30984 26382
rect 30800 26344 30802 26353
rect 30746 26279 30802 26288
rect 30930 26344 30932 26353
rect 30984 26344 30986 26353
rect 31312 26314 31340 26862
rect 30930 26279 30986 26288
rect 31300 26308 31352 26314
rect 31300 26250 31352 26256
rect 31208 26240 31260 26246
rect 31208 26182 31260 26188
rect 31220 25906 31248 26182
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 31208 25900 31260 25906
rect 31208 25842 31260 25848
rect 31024 25696 31076 25702
rect 31024 25638 31076 25644
rect 30484 22066 30604 22094
rect 30484 20534 30512 22066
rect 30472 20528 30524 20534
rect 30472 20470 30524 20476
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30392 18290 30420 19314
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30392 18034 30420 18226
rect 30300 18006 30420 18034
rect 30300 16658 30328 18006
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30484 16574 30512 20470
rect 31036 17746 31064 25638
rect 31404 22094 31432 39494
rect 31484 39432 31536 39438
rect 31484 39374 31536 39380
rect 31760 39432 31812 39438
rect 31760 39374 31812 39380
rect 31496 39098 31524 39374
rect 31484 39092 31536 39098
rect 31484 39034 31536 39040
rect 31496 38282 31524 39034
rect 31772 39030 31800 39374
rect 31760 39024 31812 39030
rect 31760 38966 31812 38972
rect 31484 38276 31536 38282
rect 31484 38218 31536 38224
rect 31864 37262 31892 39782
rect 31484 37256 31536 37262
rect 31484 37198 31536 37204
rect 31852 37256 31904 37262
rect 31852 37198 31904 37204
rect 31496 36394 31524 37198
rect 31668 37188 31720 37194
rect 31668 37130 31720 37136
rect 31680 36922 31708 37130
rect 31852 37120 31904 37126
rect 31852 37062 31904 37068
rect 31864 36922 31892 37062
rect 31668 36916 31720 36922
rect 31668 36858 31720 36864
rect 31852 36916 31904 36922
rect 31852 36858 31904 36864
rect 31496 36378 31616 36394
rect 31496 36372 31628 36378
rect 31496 36366 31576 36372
rect 31496 35630 31524 36366
rect 31576 36314 31628 36320
rect 31956 35766 31984 41414
rect 31944 35760 31996 35766
rect 31944 35702 31996 35708
rect 31852 35692 31904 35698
rect 31852 35634 31904 35640
rect 31484 35624 31536 35630
rect 31484 35566 31536 35572
rect 31496 34542 31524 35566
rect 31864 34746 31892 35634
rect 31944 35012 31996 35018
rect 31944 34954 31996 34960
rect 31852 34740 31904 34746
rect 31852 34682 31904 34688
rect 31484 34536 31536 34542
rect 31484 34478 31536 34484
rect 31760 32224 31812 32230
rect 31760 32166 31812 32172
rect 31772 31414 31800 32166
rect 31864 31414 31892 34682
rect 31956 34474 31984 34954
rect 32048 34592 32076 42026
rect 32140 41478 32168 42350
rect 32324 41592 32352 42502
rect 32416 42294 32444 43590
rect 32404 42288 32456 42294
rect 32404 42230 32456 42236
rect 32496 42220 32548 42226
rect 32496 42162 32548 42168
rect 32404 42016 32456 42022
rect 32404 41958 32456 41964
rect 32312 41586 32364 41592
rect 32312 41528 32364 41534
rect 32128 41472 32180 41478
rect 32128 41414 32180 41420
rect 32416 41414 32444 41958
rect 32324 41386 32444 41414
rect 32324 41206 32352 41386
rect 32312 41200 32364 41206
rect 32312 41142 32364 41148
rect 32128 41132 32180 41138
rect 32128 41074 32180 41080
rect 32140 40050 32168 41074
rect 32508 40526 32536 42162
rect 32600 41682 32628 45766
rect 32692 42770 32720 47620
rect 33508 47660 33560 47666
rect 33324 47602 33376 47608
rect 33428 47620 33508 47648
rect 33428 46646 33456 47620
rect 33508 47602 33560 47608
rect 33692 47660 33744 47666
rect 33692 47602 33744 47608
rect 33506 47152 33562 47161
rect 33506 47087 33508 47096
rect 33560 47087 33562 47096
rect 33508 47058 33560 47064
rect 33600 46980 33652 46986
rect 33600 46922 33652 46928
rect 33416 46640 33468 46646
rect 33416 46582 33468 46588
rect 33428 46170 33456 46582
rect 33612 46578 33640 46922
rect 33600 46572 33652 46578
rect 33600 46514 33652 46520
rect 33704 46170 33732 47602
rect 33416 46164 33468 46170
rect 33416 46106 33468 46112
rect 33692 46164 33744 46170
rect 33692 46106 33744 46112
rect 33784 45960 33836 45966
rect 33784 45902 33836 45908
rect 33692 45892 33744 45898
rect 33692 45834 33744 45840
rect 33140 45824 33192 45830
rect 33140 45766 33192 45772
rect 33152 45558 33180 45766
rect 33140 45552 33192 45558
rect 33140 45494 33192 45500
rect 33704 45286 33732 45834
rect 33796 45626 33824 45902
rect 33784 45620 33836 45626
rect 33784 45562 33836 45568
rect 33416 45280 33468 45286
rect 33692 45280 33744 45286
rect 33468 45228 33548 45234
rect 33416 45222 33548 45228
rect 33692 45222 33744 45228
rect 33428 45206 33548 45222
rect 33520 44878 33548 45206
rect 32956 44872 33008 44878
rect 32956 44814 33008 44820
rect 33508 44872 33560 44878
rect 33508 44814 33560 44820
rect 32968 44742 32996 44814
rect 32956 44736 33008 44742
rect 32956 44678 33008 44684
rect 32772 44396 32824 44402
rect 32772 44338 32824 44344
rect 32784 43926 32812 44338
rect 32772 43920 32824 43926
rect 32772 43862 32824 43868
rect 32968 43738 32996 44678
rect 33520 44402 33548 44814
rect 33508 44396 33560 44402
rect 33508 44338 33560 44344
rect 32968 43710 33088 43738
rect 32680 42764 32732 42770
rect 32680 42706 32732 42712
rect 32692 42362 32720 42706
rect 32956 42560 33008 42566
rect 32956 42502 33008 42508
rect 32680 42356 32732 42362
rect 32680 42298 32732 42304
rect 32692 41970 32720 42298
rect 32772 42016 32824 42022
rect 32692 41964 32772 41970
rect 32692 41958 32824 41964
rect 32692 41942 32812 41958
rect 32588 41676 32640 41682
rect 32588 41618 32640 41624
rect 32692 41614 32720 41942
rect 32680 41608 32732 41614
rect 32680 41550 32732 41556
rect 32588 41472 32640 41478
rect 32588 41414 32640 41420
rect 32600 41138 32628 41414
rect 32588 41132 32640 41138
rect 32588 41074 32640 41080
rect 32496 40520 32548 40526
rect 32496 40462 32548 40468
rect 32128 40044 32180 40050
rect 32128 39986 32180 39992
rect 32312 40044 32364 40050
rect 32312 39986 32364 39992
rect 32128 39568 32180 39574
rect 32128 39510 32180 39516
rect 32140 39438 32168 39510
rect 32128 39432 32180 39438
rect 32128 39374 32180 39380
rect 32220 39296 32272 39302
rect 32220 39238 32272 39244
rect 32128 37120 32180 37126
rect 32128 37062 32180 37068
rect 32140 36106 32168 37062
rect 32232 36922 32260 39238
rect 32324 39030 32352 39986
rect 32508 39438 32536 40462
rect 32600 40458 32628 41074
rect 32680 40520 32732 40526
rect 32680 40462 32732 40468
rect 32588 40452 32640 40458
rect 32588 40394 32640 40400
rect 32600 39846 32628 40394
rect 32588 39840 32640 39846
rect 32588 39782 32640 39788
rect 32496 39432 32548 39438
rect 32496 39374 32548 39380
rect 32588 39364 32640 39370
rect 32692 39352 32720 40462
rect 32772 40044 32824 40050
rect 32772 39986 32824 39992
rect 32784 39438 32812 39986
rect 32772 39432 32824 39438
rect 32772 39374 32824 39380
rect 32640 39324 32720 39352
rect 32588 39306 32640 39312
rect 32404 39296 32456 39302
rect 32404 39238 32456 39244
rect 32312 39024 32364 39030
rect 32312 38966 32364 38972
rect 32312 37324 32364 37330
rect 32312 37266 32364 37272
rect 32220 36916 32272 36922
rect 32220 36858 32272 36864
rect 32324 36666 32352 37266
rect 32416 36786 32444 39238
rect 32692 39030 32720 39324
rect 32680 39024 32732 39030
rect 32680 38966 32732 38972
rect 32496 38956 32548 38962
rect 32496 38898 32548 38904
rect 32508 38826 32536 38898
rect 32496 38820 32548 38826
rect 32496 38762 32548 38768
rect 32968 38010 32996 42502
rect 33060 41478 33088 43710
rect 33416 42900 33468 42906
rect 33416 42842 33468 42848
rect 33048 41472 33100 41478
rect 33048 41414 33100 41420
rect 33428 41138 33456 42842
rect 33508 42152 33560 42158
rect 33508 42094 33560 42100
rect 33520 41274 33548 42094
rect 33600 41744 33652 41750
rect 33600 41686 33652 41692
rect 33612 41274 33640 41686
rect 33508 41268 33560 41274
rect 33508 41210 33560 41216
rect 33600 41268 33652 41274
rect 33600 41210 33652 41216
rect 33140 41132 33192 41138
rect 33140 41074 33192 41080
rect 33416 41132 33468 41138
rect 33416 41074 33468 41080
rect 33152 40594 33180 41074
rect 33140 40588 33192 40594
rect 33140 40530 33192 40536
rect 33140 40384 33192 40390
rect 33140 40326 33192 40332
rect 33048 40044 33100 40050
rect 33048 39986 33100 39992
rect 33060 39642 33088 39986
rect 33152 39982 33180 40326
rect 33140 39976 33192 39982
rect 33140 39918 33192 39924
rect 33232 39976 33284 39982
rect 33284 39936 33364 39964
rect 33232 39918 33284 39924
rect 33048 39636 33100 39642
rect 33048 39578 33100 39584
rect 33152 39438 33180 39918
rect 33232 39840 33284 39846
rect 33232 39782 33284 39788
rect 33140 39432 33192 39438
rect 33140 39374 33192 39380
rect 33048 39092 33100 39098
rect 33048 39034 33100 39040
rect 32588 38004 32640 38010
rect 32588 37946 32640 37952
rect 32956 38004 33008 38010
rect 32956 37946 33008 37952
rect 32600 37806 32628 37946
rect 32588 37800 32640 37806
rect 32588 37742 32640 37748
rect 32956 36916 33008 36922
rect 32956 36858 33008 36864
rect 32404 36780 32456 36786
rect 32404 36722 32456 36728
rect 32324 36638 32444 36666
rect 32128 36100 32180 36106
rect 32128 36042 32180 36048
rect 32416 36038 32444 36638
rect 32864 36644 32916 36650
rect 32864 36586 32916 36592
rect 32876 36174 32904 36586
rect 32864 36168 32916 36174
rect 32864 36110 32916 36116
rect 32404 36032 32456 36038
rect 32404 35974 32456 35980
rect 32312 34604 32364 34610
rect 32048 34564 32312 34592
rect 32312 34546 32364 34552
rect 32416 34490 32444 35974
rect 32876 35766 32904 36110
rect 32864 35760 32916 35766
rect 32864 35702 32916 35708
rect 32968 35630 32996 36858
rect 32956 35624 33008 35630
rect 32956 35566 33008 35572
rect 33060 35562 33088 39034
rect 33140 37800 33192 37806
rect 33140 37742 33192 37748
rect 33152 36922 33180 37742
rect 33140 36916 33192 36922
rect 33140 36858 33192 36864
rect 33244 36106 33272 39782
rect 33336 39438 33364 39936
rect 33324 39432 33376 39438
rect 33324 39374 33376 39380
rect 33336 39302 33364 39374
rect 33324 39296 33376 39302
rect 33324 39238 33376 39244
rect 33336 38962 33364 39238
rect 33324 38956 33376 38962
rect 33324 38898 33376 38904
rect 33428 38865 33456 41074
rect 33612 40526 33640 41210
rect 33600 40520 33652 40526
rect 33600 40462 33652 40468
rect 33704 39574 33732 45222
rect 33888 40662 33916 47738
rect 34164 47666 34192 48078
rect 34152 47660 34204 47666
rect 34152 47602 34204 47608
rect 34336 44736 34388 44742
rect 34336 44678 34388 44684
rect 34150 41848 34206 41857
rect 34150 41783 34206 41792
rect 34164 41138 34192 41783
rect 34152 41132 34204 41138
rect 34152 41074 34204 41080
rect 33876 40656 33928 40662
rect 33876 40598 33928 40604
rect 33888 40390 33916 40598
rect 33876 40384 33928 40390
rect 33876 40326 33928 40332
rect 33692 39568 33744 39574
rect 33692 39510 33744 39516
rect 34348 39370 34376 44678
rect 34336 39364 34388 39370
rect 34336 39306 34388 39312
rect 33508 39296 33560 39302
rect 33508 39238 33560 39244
rect 33414 38856 33470 38865
rect 33414 38791 33470 38800
rect 33324 38344 33376 38350
rect 33324 38286 33376 38292
rect 33336 37806 33364 38286
rect 33324 37800 33376 37806
rect 33324 37742 33376 37748
rect 33416 37324 33468 37330
rect 33416 37266 33468 37272
rect 33428 36786 33456 37266
rect 33416 36780 33468 36786
rect 33416 36722 33468 36728
rect 33520 36582 33548 39238
rect 33784 38956 33836 38962
rect 33784 38898 33836 38904
rect 33600 38820 33652 38826
rect 33600 38762 33652 38768
rect 33612 38729 33640 38762
rect 33598 38720 33654 38729
rect 33598 38655 33654 38664
rect 33796 37738 33824 38898
rect 34152 38888 34204 38894
rect 34152 38830 34204 38836
rect 34242 38856 34298 38865
rect 34164 38350 34192 38830
rect 34242 38791 34244 38800
rect 34296 38791 34298 38800
rect 34244 38762 34296 38768
rect 34336 38752 34388 38758
rect 34336 38694 34388 38700
rect 34152 38344 34204 38350
rect 34348 38321 34376 38694
rect 34440 38400 34468 54538
rect 34934 53884 35242 53904
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53808 35242 53828
rect 34934 52796 35242 52816
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52720 35242 52740
rect 34934 51708 35242 51728
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51632 35242 51652
rect 34934 50620 35242 50640
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50544 35242 50564
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 35072 47184 35124 47190
rect 35072 47126 35124 47132
rect 35084 47054 35112 47126
rect 35072 47048 35124 47054
rect 35072 46990 35124 46996
rect 34704 46912 34756 46918
rect 34704 46854 34756 46860
rect 34716 46578 34744 46854
rect 35360 46646 35388 55694
rect 36740 55690 36768 59200
rect 40040 56840 40092 56846
rect 40040 56782 40092 56788
rect 40052 56438 40080 56782
rect 40040 56432 40092 56438
rect 40040 56374 40092 56380
rect 40604 56302 40632 59200
rect 42248 56840 42300 56846
rect 42248 56782 42300 56788
rect 42892 56840 42944 56846
rect 42892 56782 42944 56788
rect 40132 56296 40184 56302
rect 40132 56238 40184 56244
rect 40592 56296 40644 56302
rect 40592 56238 40644 56244
rect 40144 55894 40172 56238
rect 40132 55888 40184 55894
rect 40132 55830 40184 55836
rect 42260 55826 42288 56782
rect 42904 56438 42932 56782
rect 42892 56432 42944 56438
rect 42892 56374 42944 56380
rect 42800 56296 42852 56302
rect 42800 56238 42852 56244
rect 42248 55820 42300 55826
rect 42248 55762 42300 55768
rect 40040 55752 40092 55758
rect 40040 55694 40092 55700
rect 36268 55684 36320 55690
rect 36268 55626 36320 55632
rect 36728 55684 36780 55690
rect 36728 55626 36780 55632
rect 36280 55418 36308 55626
rect 40052 55418 40080 55694
rect 42616 55684 42668 55690
rect 42616 55626 42668 55632
rect 42628 55457 42656 55626
rect 42812 55622 42840 56238
rect 43824 55826 43852 59200
rect 44468 56438 44496 59200
rect 46664 56908 46716 56914
rect 46664 56850 46716 56856
rect 46204 56840 46256 56846
rect 46204 56782 46256 56788
rect 44456 56432 44508 56438
rect 44456 56374 44508 56380
rect 46216 55826 46244 56782
rect 46676 56370 46704 56850
rect 46664 56364 46716 56370
rect 46664 56306 46716 56312
rect 46388 56160 46440 56166
rect 46388 56102 46440 56108
rect 46400 55826 46428 56102
rect 47044 55826 47072 59200
rect 47860 56500 47912 56506
rect 47860 56442 47912 56448
rect 43812 55820 43864 55826
rect 43812 55762 43864 55768
rect 46204 55820 46256 55826
rect 46204 55762 46256 55768
rect 46388 55820 46440 55826
rect 46388 55762 46440 55768
rect 47032 55820 47084 55826
rect 47032 55762 47084 55768
rect 47872 55758 47900 56442
rect 47860 55752 47912 55758
rect 47860 55694 47912 55700
rect 42800 55616 42852 55622
rect 42800 55558 42852 55564
rect 42614 55448 42670 55457
rect 36268 55412 36320 55418
rect 36268 55354 36320 55360
rect 40040 55412 40092 55418
rect 42614 55383 42670 55392
rect 40040 55354 40092 55360
rect 36176 55276 36228 55282
rect 36176 55218 36228 55224
rect 36188 51406 36216 55218
rect 36176 51400 36228 51406
rect 36176 51342 36228 51348
rect 36084 49088 36136 49094
rect 36084 49030 36136 49036
rect 36096 48890 36124 49030
rect 36084 48884 36136 48890
rect 36084 48826 36136 48832
rect 35440 47524 35492 47530
rect 35440 47466 35492 47472
rect 35452 47122 35480 47466
rect 35532 47456 35584 47462
rect 35532 47398 35584 47404
rect 35440 47116 35492 47122
rect 35440 47058 35492 47064
rect 35544 46986 35572 47398
rect 35900 47048 35952 47054
rect 35900 46990 35952 46996
rect 35532 46980 35584 46986
rect 35532 46922 35584 46928
rect 35348 46640 35400 46646
rect 35348 46582 35400 46588
rect 34704 46572 34756 46578
rect 34704 46514 34756 46520
rect 34716 45948 34744 46514
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34888 45960 34940 45966
rect 34716 45920 34888 45948
rect 34888 45902 34940 45908
rect 34900 45490 34928 45902
rect 34888 45484 34940 45490
rect 34888 45426 34940 45432
rect 34612 45416 34664 45422
rect 34612 45358 34664 45364
rect 34624 44946 34652 45358
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34612 44940 34664 44946
rect 34612 44882 34664 44888
rect 34520 44192 34572 44198
rect 34520 44134 34572 44140
rect 34532 40118 34560 44134
rect 34624 43654 34652 44882
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34612 43648 34664 43654
rect 34612 43590 34664 43596
rect 34624 43314 34652 43590
rect 34612 43308 34664 43314
rect 34612 43250 34664 43256
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34704 42696 34756 42702
rect 34704 42638 34756 42644
rect 34716 42294 34744 42638
rect 34704 42288 34756 42294
rect 34704 42230 34756 42236
rect 34520 40112 34572 40118
rect 34520 40054 34572 40060
rect 34520 39840 34572 39846
rect 34520 39782 34572 39788
rect 34532 38457 34560 39782
rect 34612 39296 34664 39302
rect 34612 39238 34664 39244
rect 34624 38729 34652 39238
rect 34610 38720 34666 38729
rect 34610 38655 34666 38664
rect 34431 38372 34468 38400
rect 34518 38448 34574 38457
rect 34518 38383 34574 38392
rect 34152 38286 34204 38292
rect 34334 38312 34390 38321
rect 34164 37874 34192 38286
rect 34334 38247 34390 38256
rect 34336 38208 34388 38214
rect 34431 38196 34459 38372
rect 34518 38312 34574 38321
rect 34518 38247 34574 38256
rect 34431 38168 34468 38196
rect 34336 38150 34388 38156
rect 34152 37868 34204 37874
rect 34152 37810 34204 37816
rect 34164 37754 34192 37810
rect 33784 37732 33836 37738
rect 34164 37726 34284 37754
rect 33784 37674 33836 37680
rect 33796 37398 33824 37674
rect 34060 37664 34112 37670
rect 34060 37606 34112 37612
rect 34152 37664 34204 37670
rect 34152 37606 34204 37612
rect 33784 37392 33836 37398
rect 33784 37334 33836 37340
rect 33796 36786 33824 37334
rect 33968 37188 34020 37194
rect 33968 37130 34020 37136
rect 33784 36780 33836 36786
rect 33784 36722 33836 36728
rect 33980 36650 34008 37130
rect 33968 36644 34020 36650
rect 33968 36586 34020 36592
rect 33508 36576 33560 36582
rect 33508 36518 33560 36524
rect 33876 36304 33928 36310
rect 33980 36292 34008 36586
rect 33928 36264 34008 36292
rect 33876 36246 33928 36252
rect 33980 36174 34008 36264
rect 33968 36168 34020 36174
rect 33968 36110 34020 36116
rect 33232 36100 33284 36106
rect 33232 36042 33284 36048
rect 33980 35698 34008 36110
rect 33968 35692 34020 35698
rect 33968 35634 34020 35640
rect 33048 35556 33100 35562
rect 33048 35498 33100 35504
rect 33232 35488 33284 35494
rect 33232 35430 33284 35436
rect 32588 35284 32640 35290
rect 32588 35226 32640 35232
rect 32600 34610 32628 35226
rect 33244 34610 33272 35430
rect 32588 34604 32640 34610
rect 32588 34546 32640 34552
rect 33232 34604 33284 34610
rect 33232 34546 33284 34552
rect 31944 34468 31996 34474
rect 31944 34410 31996 34416
rect 32232 34462 32444 34490
rect 31760 31408 31812 31414
rect 31760 31350 31812 31356
rect 31852 31408 31904 31414
rect 31852 31350 31904 31356
rect 32232 31346 32260 34462
rect 32312 32428 32364 32434
rect 32312 32370 32364 32376
rect 32220 31340 32272 31346
rect 32220 31282 32272 31288
rect 32324 31142 32352 32370
rect 33784 31884 33836 31890
rect 33784 31826 33836 31832
rect 32496 31680 32548 31686
rect 32496 31622 32548 31628
rect 32508 31346 32536 31622
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32312 31136 32364 31142
rect 32312 31078 32364 31084
rect 31944 30184 31996 30190
rect 31944 30126 31996 30132
rect 31668 30116 31720 30122
rect 31668 30058 31720 30064
rect 31680 28994 31708 30058
rect 31852 29844 31904 29850
rect 31852 29786 31904 29792
rect 31760 29572 31812 29578
rect 31760 29514 31812 29520
rect 31772 29102 31800 29514
rect 31760 29096 31812 29102
rect 31760 29038 31812 29044
rect 31680 28966 31800 28994
rect 31484 28960 31536 28966
rect 31484 28902 31536 28908
rect 31496 28082 31524 28902
rect 31576 28212 31628 28218
rect 31576 28154 31628 28160
rect 31588 28082 31616 28154
rect 31484 28076 31536 28082
rect 31484 28018 31536 28024
rect 31576 28076 31628 28082
rect 31576 28018 31628 28024
rect 31496 27470 31524 28018
rect 31574 27840 31630 27849
rect 31574 27775 31630 27784
rect 31588 27606 31616 27775
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31576 27600 31628 27606
rect 31576 27542 31628 27548
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31576 27464 31628 27470
rect 31680 27452 31708 27610
rect 31772 27606 31800 28966
rect 31864 27674 31892 29786
rect 31956 29714 31984 30126
rect 31944 29708 31996 29714
rect 31944 29650 31996 29656
rect 32508 29578 32536 31282
rect 33796 30258 33824 31826
rect 34072 31754 34100 37606
rect 34164 37466 34192 37606
rect 34152 37460 34204 37466
rect 34152 37402 34204 37408
rect 34152 36848 34204 36854
rect 34152 36790 34204 36796
rect 34256 36802 34284 37726
rect 34348 37466 34376 38150
rect 34336 37460 34388 37466
rect 34336 37402 34388 37408
rect 34164 36378 34192 36790
rect 34256 36774 34376 36802
rect 34348 36718 34376 36774
rect 34336 36712 34388 36718
rect 34336 36654 34388 36660
rect 34152 36372 34204 36378
rect 34152 36314 34204 36320
rect 34152 35488 34204 35494
rect 34152 35430 34204 35436
rect 34164 34610 34192 35430
rect 34152 34604 34204 34610
rect 34152 34546 34204 34552
rect 34072 31726 34192 31754
rect 34164 30326 34192 31726
rect 34152 30320 34204 30326
rect 34152 30262 34204 30268
rect 33784 30252 33836 30258
rect 33784 30194 33836 30200
rect 33140 29640 33192 29646
rect 33140 29582 33192 29588
rect 33690 29608 33746 29617
rect 32496 29572 32548 29578
rect 32496 29514 32548 29520
rect 31944 29504 31996 29510
rect 31944 29446 31996 29452
rect 31956 28626 31984 29446
rect 32220 29096 32272 29102
rect 32220 29038 32272 29044
rect 31944 28620 31996 28626
rect 31944 28562 31996 28568
rect 32232 28014 32260 29038
rect 32312 28960 32364 28966
rect 32312 28902 32364 28908
rect 32324 28694 32352 28902
rect 32312 28688 32364 28694
rect 32312 28630 32364 28636
rect 32680 28552 32732 28558
rect 32680 28494 32732 28500
rect 32864 28552 32916 28558
rect 32864 28494 32916 28500
rect 32692 28218 32720 28494
rect 32680 28212 32732 28218
rect 32680 28154 32732 28160
rect 32220 28008 32272 28014
rect 32220 27950 32272 27956
rect 32680 28008 32732 28014
rect 32680 27950 32732 27956
rect 32128 27872 32180 27878
rect 32126 27840 32128 27849
rect 32180 27840 32182 27849
rect 32182 27798 32260 27826
rect 32126 27775 32182 27784
rect 31852 27668 31904 27674
rect 31852 27610 31904 27616
rect 31760 27600 31812 27606
rect 31760 27542 31812 27548
rect 31628 27424 31708 27452
rect 31576 27406 31628 27412
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31496 25906 31524 27066
rect 31668 26376 31720 26382
rect 31772 26364 31800 27542
rect 32036 27532 32088 27538
rect 31864 27492 32036 27520
rect 31864 26382 31892 27492
rect 32036 27474 32088 27480
rect 31944 27396 31996 27402
rect 31944 27338 31996 27344
rect 31720 26336 31800 26364
rect 31852 26376 31904 26382
rect 31850 26344 31852 26353
rect 31904 26344 31906 26353
rect 31668 26318 31720 26324
rect 31956 26314 31984 27338
rect 32128 27328 32180 27334
rect 32128 27270 32180 27276
rect 32140 27062 32168 27270
rect 32128 27056 32180 27062
rect 32128 26998 32180 27004
rect 32140 26518 32168 26998
rect 32232 26858 32260 27798
rect 32692 27418 32720 27950
rect 32876 27606 32904 28494
rect 33152 28422 33180 29582
rect 33690 29543 33692 29552
rect 33744 29543 33746 29552
rect 33692 29514 33744 29520
rect 33506 29064 33562 29073
rect 33506 28999 33508 29008
rect 33560 28999 33562 29008
rect 33508 28970 33560 28976
rect 33140 28416 33192 28422
rect 33140 28358 33192 28364
rect 33508 28416 33560 28422
rect 33508 28358 33560 28364
rect 33048 28076 33100 28082
rect 33048 28018 33100 28024
rect 33060 27674 33088 28018
rect 33048 27668 33100 27674
rect 33048 27610 33100 27616
rect 32864 27600 32916 27606
rect 32862 27568 32864 27577
rect 32916 27568 32918 27577
rect 32862 27503 32918 27512
rect 32496 27396 32548 27402
rect 32692 27390 32904 27418
rect 32496 27338 32548 27344
rect 32508 26926 32536 27338
rect 32876 27334 32904 27390
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 32496 26920 32548 26926
rect 32496 26862 32548 26868
rect 32220 26852 32272 26858
rect 32220 26794 32272 26800
rect 32036 26512 32088 26518
rect 32036 26454 32088 26460
rect 32128 26512 32180 26518
rect 32128 26454 32180 26460
rect 31850 26279 31906 26288
rect 31944 26308 31996 26314
rect 31944 26250 31996 26256
rect 31484 25900 31536 25906
rect 31484 25842 31536 25848
rect 32048 24274 32076 26454
rect 32232 26382 32260 26794
rect 32220 26376 32272 26382
rect 32220 26318 32272 26324
rect 32876 25838 32904 27270
rect 32864 25832 32916 25838
rect 32864 25774 32916 25780
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 32588 24132 32640 24138
rect 32588 24074 32640 24080
rect 32600 23866 32628 24074
rect 32588 23860 32640 23866
rect 32588 23802 32640 23808
rect 33152 23730 33180 28358
rect 33520 28150 33548 28358
rect 33508 28144 33560 28150
rect 33508 28086 33560 28092
rect 33796 28082 33824 30194
rect 34058 28248 34114 28257
rect 34058 28183 34114 28192
rect 34072 28150 34100 28183
rect 34060 28144 34112 28150
rect 34060 28086 34112 28092
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 34440 27878 34468 38168
rect 34532 36378 34560 38247
rect 34612 38208 34664 38214
rect 34612 38150 34664 38156
rect 34520 36372 34572 36378
rect 34520 36314 34572 36320
rect 34520 36168 34572 36174
rect 34520 36110 34572 36116
rect 34532 31822 34560 36110
rect 34624 33998 34652 38150
rect 34716 36242 34744 42230
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34888 40656 34940 40662
rect 34888 40598 34940 40604
rect 34796 40384 34848 40390
rect 34796 40326 34848 40332
rect 34808 39506 34836 40326
rect 34900 39982 34928 40598
rect 34980 40452 35032 40458
rect 34980 40394 35032 40400
rect 34992 39982 35020 40394
rect 34888 39976 34940 39982
rect 34888 39918 34940 39924
rect 34980 39976 35032 39982
rect 34980 39918 35032 39924
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34796 39500 34848 39506
rect 34796 39442 34848 39448
rect 34888 39432 34940 39438
rect 34888 39374 34940 39380
rect 34900 38962 34928 39374
rect 34888 38956 34940 38962
rect 34888 38898 34940 38904
rect 34796 38752 34848 38758
rect 34796 38694 34848 38700
rect 34808 38554 34836 38694
rect 35360 38677 35388 46582
rect 35912 46510 35940 46990
rect 36188 46714 36216 51342
rect 37832 49836 37884 49842
rect 37832 49778 37884 49784
rect 39212 49836 39264 49842
rect 39212 49778 39264 49784
rect 39948 49836 40000 49842
rect 39948 49778 40000 49784
rect 40316 49836 40368 49842
rect 40316 49778 40368 49784
rect 37372 49768 37424 49774
rect 37372 49710 37424 49716
rect 37384 49230 37412 49710
rect 37372 49224 37424 49230
rect 37372 49166 37424 49172
rect 37280 49156 37332 49162
rect 37280 49098 37332 49104
rect 37292 48346 37320 49098
rect 37384 48754 37412 49166
rect 37372 48748 37424 48754
rect 37372 48690 37424 48696
rect 37280 48340 37332 48346
rect 37280 48282 37332 48288
rect 36544 48136 36596 48142
rect 37188 48136 37240 48142
rect 36544 48078 36596 48084
rect 37108 48096 37188 48124
rect 36176 46708 36228 46714
rect 36176 46650 36228 46656
rect 35900 46504 35952 46510
rect 35900 46446 35952 46452
rect 35808 46096 35860 46102
rect 35808 46038 35860 46044
rect 35532 45824 35584 45830
rect 35532 45766 35584 45772
rect 35544 45472 35572 45766
rect 35624 45484 35676 45490
rect 35544 45444 35624 45472
rect 35440 45280 35492 45286
rect 35440 45222 35492 45228
rect 35452 45082 35480 45222
rect 35440 45076 35492 45082
rect 35440 45018 35492 45024
rect 35544 44402 35572 45444
rect 35624 45426 35676 45432
rect 35624 45348 35676 45354
rect 35624 45290 35676 45296
rect 35636 44742 35664 45290
rect 35716 45280 35768 45286
rect 35716 45222 35768 45228
rect 35728 44878 35756 45222
rect 35716 44872 35768 44878
rect 35716 44814 35768 44820
rect 35624 44736 35676 44742
rect 35624 44678 35676 44684
rect 35820 44402 35848 46038
rect 35532 44396 35584 44402
rect 35532 44338 35584 44344
rect 35808 44396 35860 44402
rect 35808 44338 35860 44344
rect 35544 43994 35572 44338
rect 35532 43988 35584 43994
rect 35532 43930 35584 43936
rect 35544 43314 35572 43930
rect 35912 43790 35940 46446
rect 35992 45960 36044 45966
rect 35992 45902 36044 45908
rect 36004 45286 36032 45902
rect 36268 45824 36320 45830
rect 36268 45766 36320 45772
rect 35992 45280 36044 45286
rect 35992 45222 36044 45228
rect 35990 44432 36046 44441
rect 35990 44367 35992 44376
rect 36044 44367 36046 44376
rect 35992 44338 36044 44344
rect 35900 43784 35952 43790
rect 35900 43726 35952 43732
rect 35532 43308 35584 43314
rect 35532 43250 35584 43256
rect 35624 43240 35676 43246
rect 35624 43182 35676 43188
rect 35440 43172 35492 43178
rect 35440 43114 35492 43120
rect 35452 40202 35480 43114
rect 35532 43104 35584 43110
rect 35532 43046 35584 43052
rect 35544 42226 35572 43046
rect 35636 42362 35664 43182
rect 35912 42838 35940 43726
rect 35992 43648 36044 43654
rect 35992 43590 36044 43596
rect 36004 43314 36032 43590
rect 36280 43314 36308 45766
rect 36452 45484 36504 45490
rect 36452 45426 36504 45432
rect 36464 45393 36492 45426
rect 36450 45384 36506 45393
rect 36450 45319 36506 45328
rect 36452 45280 36504 45286
rect 36450 45248 36452 45257
rect 36504 45248 36506 45257
rect 36450 45183 36506 45192
rect 35992 43308 36044 43314
rect 35992 43250 36044 43256
rect 36268 43308 36320 43314
rect 36268 43250 36320 43256
rect 36084 43240 36136 43246
rect 36084 43182 36136 43188
rect 35900 42832 35952 42838
rect 35900 42774 35952 42780
rect 36096 42566 36124 43182
rect 36084 42560 36136 42566
rect 36084 42502 36136 42508
rect 35624 42356 35676 42362
rect 35624 42298 35676 42304
rect 35532 42220 35584 42226
rect 35532 42162 35584 42168
rect 35636 41206 35664 42298
rect 35624 41200 35676 41206
rect 35624 41142 35676 41148
rect 35452 40174 35664 40202
rect 35440 40044 35492 40050
rect 35440 39986 35492 39992
rect 35452 39574 35480 39986
rect 35440 39568 35492 39574
rect 35440 39510 35492 39516
rect 35440 39092 35492 39098
rect 35440 39034 35492 39040
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 35346 38668 35402 38677
rect 35346 38603 35402 38612
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34796 38548 34848 38554
rect 34796 38490 34848 38496
rect 35162 38448 35218 38457
rect 35162 38383 35164 38392
rect 35216 38383 35218 38392
rect 35164 38354 35216 38360
rect 35346 38312 35402 38321
rect 35346 38247 35402 38256
rect 34796 38208 34848 38214
rect 34796 38150 34848 38156
rect 34808 37330 34836 38150
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 34808 36718 34836 37062
rect 35256 36780 35308 36786
rect 35256 36722 35308 36728
rect 34796 36712 34848 36718
rect 34796 36654 34848 36660
rect 35268 36650 35296 36722
rect 35256 36644 35308 36650
rect 35256 36586 35308 36592
rect 34796 36576 34848 36582
rect 34796 36518 34848 36524
rect 34704 36236 34756 36242
rect 34704 36178 34756 36184
rect 34716 35154 34744 36178
rect 34808 36174 34836 36518
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34980 36304 35032 36310
rect 34980 36246 35032 36252
rect 34796 36168 34848 36174
rect 34796 36110 34848 36116
rect 34796 36032 34848 36038
rect 34796 35974 34848 35980
rect 34704 35148 34756 35154
rect 34704 35090 34756 35096
rect 34716 34066 34744 35090
rect 34704 34060 34756 34066
rect 34704 34002 34756 34008
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34716 32502 34744 34002
rect 34704 32496 34756 32502
rect 34704 32438 34756 32444
rect 34716 31890 34744 32438
rect 34808 32434 34836 35974
rect 34992 35766 35020 36246
rect 35256 36168 35308 36174
rect 35256 36110 35308 36116
rect 34980 35760 35032 35766
rect 34980 35702 35032 35708
rect 35268 35698 35296 36110
rect 35256 35692 35308 35698
rect 35256 35634 35308 35640
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34796 32428 34848 32434
rect 34796 32370 34848 32376
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34704 31884 34756 31890
rect 34704 31826 34756 31832
rect 34520 31816 34572 31822
rect 34520 31758 34572 31764
rect 34716 31754 34744 31826
rect 34704 31748 34756 31754
rect 34704 31690 34756 31696
rect 34980 31680 35032 31686
rect 34980 31622 35032 31628
rect 34992 31346 35020 31622
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34980 31340 35032 31346
rect 34980 31282 35032 31288
rect 34716 30734 34744 31282
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34704 30728 34756 30734
rect 34704 30670 34756 30676
rect 34716 28626 34744 30670
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34704 28620 34756 28626
rect 34704 28562 34756 28568
rect 34428 27872 34480 27878
rect 34428 27814 34480 27820
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34152 24132 34204 24138
rect 34152 24074 34204 24080
rect 33140 23724 33192 23730
rect 33140 23666 33192 23672
rect 31128 22066 31432 22094
rect 31128 19922 31156 22066
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31116 19916 31168 19922
rect 31116 19858 31168 19864
rect 31220 19802 31248 20946
rect 31128 19774 31248 19802
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 30484 16546 30604 16574
rect 29840 6886 29960 6914
rect 29460 6316 29512 6322
rect 29460 6258 29512 6264
rect 29840 4146 29868 6886
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 29184 4072 29236 4078
rect 29184 4014 29236 4020
rect 30576 4010 30604 16546
rect 31128 4146 31156 19774
rect 31208 18080 31260 18086
rect 31208 18022 31260 18028
rect 31220 17746 31248 18022
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 32864 17604 32916 17610
rect 32864 17546 32916 17552
rect 32876 16574 32904 17546
rect 32876 16546 32996 16574
rect 31116 4140 31168 4146
rect 31116 4082 31168 4088
rect 30564 4004 30616 4010
rect 30564 3946 30616 3952
rect 29736 3936 29788 3942
rect 29736 3878 29788 3884
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 32128 3936 32180 3942
rect 32128 3878 32180 3884
rect 28816 3460 28868 3466
rect 28816 3402 28868 3408
rect 28828 2854 28856 3402
rect 29748 3058 29776 3878
rect 30668 3602 30696 3878
rect 30656 3596 30708 3602
rect 30656 3538 30708 3544
rect 30760 3126 30788 3878
rect 32140 3602 32168 3878
rect 32968 3670 32996 16546
rect 32956 3664 33008 3670
rect 32956 3606 33008 3612
rect 34164 3602 34192 24074
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35360 21010 35388 38247
rect 35452 35018 35480 39034
rect 35636 38826 35664 40174
rect 35808 39364 35860 39370
rect 35808 39306 35860 39312
rect 35716 38888 35768 38894
rect 35716 38830 35768 38836
rect 35624 38820 35676 38826
rect 35624 38762 35676 38768
rect 35532 38752 35584 38758
rect 35532 38694 35584 38700
rect 35544 35630 35572 38694
rect 35624 38344 35676 38350
rect 35624 38286 35676 38292
rect 35636 36786 35664 38286
rect 35728 37874 35756 38830
rect 35820 37942 35848 39306
rect 35992 39296 36044 39302
rect 35992 39238 36044 39244
rect 35900 38208 35952 38214
rect 35900 38150 35952 38156
rect 35808 37936 35860 37942
rect 35808 37878 35860 37884
rect 35716 37868 35768 37874
rect 35716 37810 35768 37816
rect 35728 37262 35756 37810
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35820 36854 35848 37878
rect 35808 36848 35860 36854
rect 35808 36790 35860 36796
rect 35624 36780 35676 36786
rect 35624 36722 35676 36728
rect 35716 36712 35768 36718
rect 35716 36654 35768 36660
rect 35624 36576 35676 36582
rect 35624 36518 35676 36524
rect 35532 35624 35584 35630
rect 35532 35566 35584 35572
rect 35440 35012 35492 35018
rect 35440 34954 35492 34960
rect 35532 34536 35584 34542
rect 35532 34478 35584 34484
rect 35544 30734 35572 34478
rect 35532 30728 35584 30734
rect 35532 30670 35584 30676
rect 35544 30394 35572 30670
rect 35532 30388 35584 30394
rect 35532 30330 35584 30336
rect 35636 28490 35664 36518
rect 35728 36378 35756 36654
rect 35716 36372 35768 36378
rect 35716 36314 35768 36320
rect 35820 35834 35848 36790
rect 35808 35828 35860 35834
rect 35808 35770 35860 35776
rect 35716 34672 35768 34678
rect 35716 34614 35768 34620
rect 35728 32434 35756 34614
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35716 32428 35768 32434
rect 35716 32370 35768 32376
rect 35728 31686 35756 32370
rect 35820 31754 35848 32846
rect 35808 31748 35860 31754
rect 35808 31690 35860 31696
rect 35716 31680 35768 31686
rect 35716 31622 35768 31628
rect 35820 31346 35848 31690
rect 35912 31482 35940 38150
rect 36004 36650 36032 39238
rect 36096 39030 36124 42502
rect 36084 39024 36136 39030
rect 36084 38966 36136 38972
rect 36556 38418 36584 48078
rect 36728 46368 36780 46374
rect 36728 46310 36780 46316
rect 36636 45824 36688 45830
rect 36636 45766 36688 45772
rect 36648 45490 36676 45766
rect 36740 45490 36768 46310
rect 37004 45960 37056 45966
rect 37004 45902 37056 45908
rect 36636 45484 36688 45490
rect 36636 45426 36688 45432
rect 36728 45484 36780 45490
rect 36728 45426 36780 45432
rect 37016 45286 37044 45902
rect 37004 45280 37056 45286
rect 37004 45222 37056 45228
rect 36728 43104 36780 43110
rect 36728 43046 36780 43052
rect 36740 42702 36768 43046
rect 36728 42696 36780 42702
rect 36728 42638 36780 42644
rect 36820 39976 36872 39982
rect 36820 39918 36872 39924
rect 36728 38548 36780 38554
rect 36728 38490 36780 38496
rect 36544 38412 36596 38418
rect 36544 38354 36596 38360
rect 36268 38344 36320 38350
rect 36268 38286 36320 38292
rect 36636 38344 36688 38350
rect 36636 38286 36688 38292
rect 36280 38010 36308 38286
rect 36268 38004 36320 38010
rect 36268 37946 36320 37952
rect 36648 37942 36676 38286
rect 36740 38282 36768 38490
rect 36728 38276 36780 38282
rect 36728 38218 36780 38224
rect 36636 37936 36688 37942
rect 36636 37878 36688 37884
rect 36176 37868 36228 37874
rect 36176 37810 36228 37816
rect 36452 37868 36504 37874
rect 36452 37810 36504 37816
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 35992 36644 36044 36650
rect 35992 36586 36044 36592
rect 36096 36242 36124 37198
rect 36188 37126 36216 37810
rect 36464 37466 36492 37810
rect 36728 37664 36780 37670
rect 36728 37606 36780 37612
rect 36452 37460 36504 37466
rect 36452 37402 36504 37408
rect 36360 37324 36412 37330
rect 36360 37266 36412 37272
rect 36176 37120 36228 37126
rect 36176 37062 36228 37068
rect 36372 36854 36400 37266
rect 36360 36848 36412 36854
rect 36360 36790 36412 36796
rect 36542 36816 36598 36825
rect 36176 36780 36228 36786
rect 36176 36722 36228 36728
rect 36452 36780 36504 36786
rect 36542 36751 36544 36760
rect 36452 36722 36504 36728
rect 36596 36751 36598 36760
rect 36544 36722 36596 36728
rect 36084 36236 36136 36242
rect 36084 36178 36136 36184
rect 35992 36100 36044 36106
rect 35992 36042 36044 36048
rect 36004 35494 36032 36042
rect 36188 35562 36216 36722
rect 36464 36378 36492 36722
rect 36452 36372 36504 36378
rect 36452 36314 36504 36320
rect 36176 35556 36228 35562
rect 36176 35498 36228 35504
rect 35992 35488 36044 35494
rect 35992 35430 36044 35436
rect 36082 33960 36138 33969
rect 36082 33895 36138 33904
rect 36096 33862 36124 33895
rect 36084 33856 36136 33862
rect 36084 33798 36136 33804
rect 36740 32502 36768 37606
rect 36832 36174 36860 39918
rect 37108 38865 37136 48096
rect 37188 48078 37240 48084
rect 37372 48000 37424 48006
rect 37372 47942 37424 47948
rect 37384 47666 37412 47942
rect 37844 47802 37872 49778
rect 38936 49632 38988 49638
rect 38936 49574 38988 49580
rect 38948 49298 38976 49574
rect 38936 49292 38988 49298
rect 38936 49234 38988 49240
rect 38752 49088 38804 49094
rect 38752 49030 38804 49036
rect 38764 48754 38792 49030
rect 38200 48748 38252 48754
rect 38200 48690 38252 48696
rect 38752 48748 38804 48754
rect 38752 48690 38804 48696
rect 38212 48346 38240 48690
rect 39224 48686 39252 49778
rect 39672 49768 39724 49774
rect 39672 49710 39724 49716
rect 39212 48680 39264 48686
rect 39212 48622 39264 48628
rect 38200 48340 38252 48346
rect 38200 48282 38252 48288
rect 38108 48136 38160 48142
rect 38108 48078 38160 48084
rect 37832 47796 37884 47802
rect 37832 47738 37884 47744
rect 37556 47728 37608 47734
rect 37556 47670 37608 47676
rect 37280 47660 37332 47666
rect 37280 47602 37332 47608
rect 37372 47660 37424 47666
rect 37372 47602 37424 47608
rect 37292 47190 37320 47602
rect 37568 47462 37596 47670
rect 38120 47666 38148 48078
rect 39224 47666 39252 48622
rect 39684 48074 39712 49710
rect 39960 49434 39988 49778
rect 39948 49428 40000 49434
rect 39948 49370 40000 49376
rect 39856 49292 39908 49298
rect 39856 49234 39908 49240
rect 39764 48272 39816 48278
rect 39764 48214 39816 48220
rect 39672 48068 39724 48074
rect 39672 48010 39724 48016
rect 38108 47660 38160 47666
rect 38108 47602 38160 47608
rect 39212 47660 39264 47666
rect 39212 47602 39264 47608
rect 37556 47456 37608 47462
rect 37556 47398 37608 47404
rect 39776 47190 39804 48214
rect 39868 47530 39896 49234
rect 40328 49230 40356 49778
rect 41512 49768 41564 49774
rect 41512 49710 41564 49716
rect 40132 49224 40184 49230
rect 40132 49166 40184 49172
rect 40316 49224 40368 49230
rect 40316 49166 40368 49172
rect 39948 48748 40000 48754
rect 39948 48690 40000 48696
rect 39960 48142 39988 48690
rect 40144 48686 40172 49166
rect 40132 48680 40184 48686
rect 40132 48622 40184 48628
rect 40592 48680 40644 48686
rect 40592 48622 40644 48628
rect 41144 48680 41196 48686
rect 41144 48622 41196 48628
rect 40604 48142 40632 48622
rect 40684 48544 40736 48550
rect 40684 48486 40736 48492
rect 39948 48136 40000 48142
rect 39948 48078 40000 48084
rect 40592 48136 40644 48142
rect 40592 48078 40644 48084
rect 40604 47734 40632 48078
rect 40592 47728 40644 47734
rect 40592 47670 40644 47676
rect 39856 47524 39908 47530
rect 39856 47466 39908 47472
rect 37280 47184 37332 47190
rect 37280 47126 37332 47132
rect 37648 47184 37700 47190
rect 37648 47126 37700 47132
rect 39764 47184 39816 47190
rect 39764 47126 39816 47132
rect 37280 46572 37332 46578
rect 37280 46514 37332 46520
rect 37188 45892 37240 45898
rect 37188 45834 37240 45840
rect 37200 45082 37228 45834
rect 37292 45234 37320 46514
rect 37292 45206 37412 45234
rect 37188 45076 37240 45082
rect 37188 45018 37240 45024
rect 37280 41608 37332 41614
rect 37280 41550 37332 41556
rect 37292 40730 37320 41550
rect 37280 40724 37332 40730
rect 37280 40666 37332 40672
rect 37188 40520 37240 40526
rect 37188 40462 37240 40468
rect 37200 40390 37228 40462
rect 37188 40384 37240 40390
rect 37188 40326 37240 40332
rect 37280 39432 37332 39438
rect 37280 39374 37332 39380
rect 37292 38962 37320 39374
rect 37384 39302 37412 45206
rect 37556 44872 37608 44878
rect 37556 44814 37608 44820
rect 37568 43994 37596 44814
rect 37556 43988 37608 43994
rect 37556 43930 37608 43936
rect 37556 42764 37608 42770
rect 37556 42706 37608 42712
rect 37568 41614 37596 42706
rect 37556 41608 37608 41614
rect 37556 41550 37608 41556
rect 37660 41414 37688 47126
rect 39776 47054 39804 47126
rect 39672 47048 39724 47054
rect 39670 47016 39672 47025
rect 39764 47048 39816 47054
rect 39724 47016 39726 47025
rect 37924 46980 37976 46986
rect 40316 47048 40368 47054
rect 39764 46990 39816 46996
rect 40144 47008 40316 47036
rect 39670 46951 39726 46960
rect 37924 46922 37976 46928
rect 37936 46578 37964 46922
rect 39304 46708 39356 46714
rect 39304 46650 39356 46656
rect 39210 46608 39266 46617
rect 37924 46572 37976 46578
rect 39210 46543 39212 46552
rect 37924 46514 37976 46520
rect 39264 46543 39266 46552
rect 39212 46514 39264 46520
rect 38844 46436 38896 46442
rect 38844 46378 38896 46384
rect 38476 46368 38528 46374
rect 38476 46310 38528 46316
rect 38384 46164 38436 46170
rect 38384 46106 38436 46112
rect 37832 45960 37884 45966
rect 37832 45902 37884 45908
rect 38108 45960 38160 45966
rect 38108 45902 38160 45908
rect 37740 45824 37792 45830
rect 37740 45766 37792 45772
rect 37752 45490 37780 45766
rect 37740 45484 37792 45490
rect 37740 45426 37792 45432
rect 37752 44946 37780 45426
rect 37740 44940 37792 44946
rect 37740 44882 37792 44888
rect 37844 44878 37872 45902
rect 37924 45824 37976 45830
rect 37924 45766 37976 45772
rect 37936 45626 37964 45766
rect 37924 45620 37976 45626
rect 37924 45562 37976 45568
rect 37922 45384 37978 45393
rect 37922 45319 37924 45328
rect 37976 45319 37978 45328
rect 38016 45348 38068 45354
rect 37924 45290 37976 45296
rect 38016 45290 38068 45296
rect 37936 44946 37964 45290
rect 38028 45082 38056 45290
rect 38120 45098 38148 45902
rect 38292 45484 38344 45490
rect 38292 45426 38344 45432
rect 38200 45280 38252 45286
rect 38198 45248 38200 45257
rect 38252 45248 38254 45257
rect 38198 45183 38254 45192
rect 38016 45076 38068 45082
rect 38120 45070 38240 45098
rect 38016 45018 38068 45024
rect 37924 44940 37976 44946
rect 37924 44882 37976 44888
rect 38212 44878 38240 45070
rect 37832 44872 37884 44878
rect 37832 44814 37884 44820
rect 38200 44872 38252 44878
rect 38200 44814 38252 44820
rect 37844 44470 37872 44814
rect 37832 44464 37884 44470
rect 37832 44406 37884 44412
rect 37740 43104 37792 43110
rect 37740 43046 37792 43052
rect 37752 42906 37780 43046
rect 37740 42900 37792 42906
rect 37740 42842 37792 42848
rect 37844 42226 37872 44406
rect 38304 44266 38332 45426
rect 38396 45082 38424 46106
rect 38488 45966 38516 46310
rect 38476 45960 38528 45966
rect 38476 45902 38528 45908
rect 38384 45076 38436 45082
rect 38384 45018 38436 45024
rect 38384 44872 38436 44878
rect 38384 44814 38436 44820
rect 38396 44334 38424 44814
rect 38488 44810 38516 45902
rect 38752 45892 38804 45898
rect 38752 45834 38804 45840
rect 38764 45626 38792 45834
rect 38752 45620 38804 45626
rect 38752 45562 38804 45568
rect 38568 45484 38620 45490
rect 38568 45426 38620 45432
rect 38476 44804 38528 44810
rect 38476 44746 38528 44752
rect 38580 44538 38608 45426
rect 38660 45280 38712 45286
rect 38660 45222 38712 45228
rect 38672 44878 38700 45222
rect 38660 44872 38712 44878
rect 38660 44814 38712 44820
rect 38568 44532 38620 44538
rect 38568 44474 38620 44480
rect 38384 44328 38436 44334
rect 38384 44270 38436 44276
rect 38292 44260 38344 44266
rect 38292 44202 38344 44208
rect 38108 43784 38160 43790
rect 38108 43726 38160 43732
rect 37832 42220 37884 42226
rect 37832 42162 37884 42168
rect 37924 41608 37976 41614
rect 37924 41550 37976 41556
rect 37568 41386 37688 41414
rect 37372 39296 37424 39302
rect 37372 39238 37424 39244
rect 37568 38978 37596 41386
rect 37936 41138 37964 41550
rect 37924 41132 37976 41138
rect 37924 41074 37976 41080
rect 37832 41064 37884 41070
rect 37832 41006 37884 41012
rect 37844 40594 37872 41006
rect 37936 40594 37964 41074
rect 37832 40588 37884 40594
rect 37832 40530 37884 40536
rect 37924 40588 37976 40594
rect 37924 40530 37976 40536
rect 37936 40186 37964 40530
rect 37924 40180 37976 40186
rect 37924 40122 37976 40128
rect 37740 39296 37792 39302
rect 37740 39238 37792 39244
rect 37648 39092 37700 39098
rect 37648 39034 37700 39040
rect 37280 38956 37332 38962
rect 37280 38898 37332 38904
rect 37384 38950 37596 38978
rect 37094 38856 37150 38865
rect 37094 38791 37150 38800
rect 37108 38654 37136 38791
rect 37108 38626 37320 38654
rect 37292 38350 37320 38626
rect 37280 38344 37332 38350
rect 37280 38286 37332 38292
rect 37096 38208 37148 38214
rect 37384 38196 37412 38950
rect 37660 38842 37688 39034
rect 37568 38814 37688 38842
rect 37568 38486 37596 38814
rect 37648 38752 37700 38758
rect 37648 38694 37700 38700
rect 37556 38480 37608 38486
rect 37556 38422 37608 38428
rect 37568 38282 37596 38422
rect 37556 38276 37608 38282
rect 37556 38218 37608 38224
rect 37096 38150 37148 38156
rect 37200 38168 37412 38196
rect 36820 36168 36872 36174
rect 36820 36110 36872 36116
rect 36728 32496 36780 32502
rect 36728 32438 36780 32444
rect 36728 32224 36780 32230
rect 36728 32166 36780 32172
rect 35900 31476 35952 31482
rect 35900 31418 35952 31424
rect 35808 31340 35860 31346
rect 35808 31282 35860 31288
rect 36636 31136 36688 31142
rect 36636 31078 36688 31084
rect 36648 30734 36676 31078
rect 36740 30938 36768 32166
rect 36728 30932 36780 30938
rect 36728 30874 36780 30880
rect 36740 30734 36768 30874
rect 36636 30728 36688 30734
rect 36636 30670 36688 30676
rect 36728 30728 36780 30734
rect 36728 30670 36780 30676
rect 35808 30048 35860 30054
rect 35808 29990 35860 29996
rect 36452 30048 36504 30054
rect 36452 29990 36504 29996
rect 35820 28626 35848 29990
rect 36464 29782 36492 29990
rect 36452 29776 36504 29782
rect 36452 29718 36504 29724
rect 36648 29714 36676 30670
rect 36636 29708 36688 29714
rect 36636 29650 36688 29656
rect 36268 29504 36320 29510
rect 36268 29446 36320 29452
rect 35808 28620 35860 28626
rect 35808 28562 35860 28568
rect 35624 28484 35676 28490
rect 35624 28426 35676 28432
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 36188 28082 36216 28358
rect 36176 28076 36228 28082
rect 36176 28018 36228 28024
rect 36188 27606 36216 28018
rect 36176 27600 36228 27606
rect 36176 27542 36228 27548
rect 36280 27452 36308 29446
rect 36728 29028 36780 29034
rect 36728 28970 36780 28976
rect 36360 28076 36412 28082
rect 36360 28018 36412 28024
rect 36372 27674 36400 28018
rect 36544 27872 36596 27878
rect 36544 27814 36596 27820
rect 36360 27668 36412 27674
rect 36360 27610 36412 27616
rect 36360 27464 36412 27470
rect 36280 27424 36360 27452
rect 36360 27406 36412 27412
rect 36556 26858 36584 27814
rect 36740 27334 36768 28970
rect 36832 28694 36860 36110
rect 37108 32910 37136 38150
rect 37200 37806 37228 38168
rect 37188 37800 37240 37806
rect 37188 37742 37240 37748
rect 37372 37800 37424 37806
rect 37372 37742 37424 37748
rect 37384 37398 37412 37742
rect 37568 37738 37596 38218
rect 37556 37732 37608 37738
rect 37556 37674 37608 37680
rect 37464 37664 37516 37670
rect 37464 37606 37516 37612
rect 37372 37392 37424 37398
rect 37372 37334 37424 37340
rect 37280 37256 37332 37262
rect 37280 37198 37332 37204
rect 37292 36310 37320 37198
rect 37384 36825 37412 37334
rect 37370 36816 37426 36825
rect 37370 36751 37372 36760
rect 37424 36751 37426 36760
rect 37372 36722 37424 36728
rect 37384 36691 37412 36722
rect 37372 36576 37424 36582
rect 37372 36518 37424 36524
rect 37280 36304 37332 36310
rect 37280 36246 37332 36252
rect 37384 35698 37412 36518
rect 37372 35692 37424 35698
rect 37372 35634 37424 35640
rect 37280 35624 37332 35630
rect 37280 35566 37332 35572
rect 37292 35086 37320 35566
rect 37280 35080 37332 35086
rect 37280 35022 37332 35028
rect 37188 34944 37240 34950
rect 37188 34886 37240 34892
rect 37200 33561 37228 34886
rect 37186 33552 37242 33561
rect 37186 33487 37242 33496
rect 37096 32904 37148 32910
rect 37096 32846 37148 32852
rect 37188 32428 37240 32434
rect 37188 32370 37240 32376
rect 37200 31890 37228 32370
rect 37188 31884 37240 31890
rect 37188 31826 37240 31832
rect 37476 31822 37504 37606
rect 37568 37330 37596 37674
rect 37556 37324 37608 37330
rect 37556 37266 37608 37272
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 37660 31414 37688 38694
rect 37752 36854 37780 39238
rect 37832 38956 37884 38962
rect 37832 38898 37884 38904
rect 37844 38350 37872 38898
rect 37832 38344 37884 38350
rect 37832 38286 37884 38292
rect 37844 37942 37872 38286
rect 37832 37936 37884 37942
rect 37832 37878 37884 37884
rect 37740 36848 37792 36854
rect 37740 36790 37792 36796
rect 37832 36576 37884 36582
rect 37832 36518 37884 36524
rect 37844 35086 37872 36518
rect 37832 35080 37884 35086
rect 37832 35022 37884 35028
rect 37648 31408 37700 31414
rect 37648 31350 37700 31356
rect 37188 30660 37240 30666
rect 37188 30602 37240 30608
rect 37096 30592 37148 30598
rect 37096 30534 37148 30540
rect 37108 30326 37136 30534
rect 37096 30320 37148 30326
rect 37096 30262 37148 30268
rect 37200 29646 37228 30602
rect 37648 30048 37700 30054
rect 37648 29990 37700 29996
rect 37740 30048 37792 30054
rect 37740 29990 37792 29996
rect 37004 29640 37056 29646
rect 37004 29582 37056 29588
rect 37188 29640 37240 29646
rect 37188 29582 37240 29588
rect 37016 29034 37044 29582
rect 37372 29096 37424 29102
rect 37372 29038 37424 29044
rect 37004 29028 37056 29034
rect 37004 28970 37056 28976
rect 36820 28688 36872 28694
rect 36820 28630 36872 28636
rect 36728 27328 36780 27334
rect 36728 27270 36780 27276
rect 36740 26994 36768 27270
rect 36832 27062 36860 28630
rect 37384 28506 37412 29038
rect 37464 28960 37516 28966
rect 37464 28902 37516 28908
rect 37292 28490 37412 28506
rect 37188 28484 37240 28490
rect 37188 28426 37240 28432
rect 37280 28484 37412 28490
rect 37332 28478 37412 28484
rect 37280 28426 37332 28432
rect 37200 27946 37228 28426
rect 37292 28082 37320 28426
rect 37476 28082 37504 28902
rect 37280 28076 37332 28082
rect 37280 28018 37332 28024
rect 37464 28076 37516 28082
rect 37464 28018 37516 28024
rect 37660 27962 37688 29990
rect 37752 28558 37780 29990
rect 37924 29164 37976 29170
rect 37924 29106 37976 29112
rect 37740 28552 37792 28558
rect 37740 28494 37792 28500
rect 37752 28150 37780 28494
rect 37740 28144 37792 28150
rect 37740 28086 37792 28092
rect 37936 28082 37964 29106
rect 38016 28960 38068 28966
rect 38016 28902 38068 28908
rect 38028 28558 38056 28902
rect 38016 28552 38068 28558
rect 38016 28494 38068 28500
rect 38120 28422 38148 43726
rect 38292 43716 38344 43722
rect 38292 43658 38344 43664
rect 38384 43716 38436 43722
rect 38384 43658 38436 43664
rect 38200 42220 38252 42226
rect 38200 42162 38252 42168
rect 38212 41274 38240 42162
rect 38200 41268 38252 41274
rect 38200 41210 38252 41216
rect 38304 31754 38332 43658
rect 38396 43314 38424 43658
rect 38384 43308 38436 43314
rect 38384 43250 38436 43256
rect 38384 42764 38436 42770
rect 38384 42706 38436 42712
rect 38396 41818 38424 42706
rect 38580 42702 38608 44474
rect 38752 43784 38804 43790
rect 38856 43772 38884 46378
rect 39316 46374 39344 46650
rect 39776 46578 39804 46990
rect 40144 46578 40172 47008
rect 40316 46990 40368 46996
rect 40316 46912 40368 46918
rect 40316 46854 40368 46860
rect 40328 46578 40356 46854
rect 39764 46572 39816 46578
rect 39764 46514 39816 46520
rect 40132 46572 40184 46578
rect 40132 46514 40184 46520
rect 40316 46572 40368 46578
rect 40316 46514 40368 46520
rect 39304 46368 39356 46374
rect 39304 46310 39356 46316
rect 39120 46028 39172 46034
rect 39120 45970 39172 45976
rect 38936 45960 38988 45966
rect 38936 45902 38988 45908
rect 38948 43994 38976 45902
rect 39132 45422 39160 45970
rect 40040 45892 40092 45898
rect 40040 45834 40092 45840
rect 39856 45824 39908 45830
rect 39856 45766 39908 45772
rect 39868 45626 39896 45766
rect 39856 45620 39908 45626
rect 39856 45562 39908 45568
rect 40052 45558 40080 45834
rect 39948 45552 40000 45558
rect 39946 45520 39948 45529
rect 40040 45552 40092 45558
rect 40000 45520 40002 45529
rect 39764 45484 39816 45490
rect 40040 45494 40092 45500
rect 39946 45455 40002 45464
rect 39764 45426 39816 45432
rect 39120 45416 39172 45422
rect 39120 45358 39172 45364
rect 39132 45082 39160 45358
rect 39120 45076 39172 45082
rect 39120 45018 39172 45024
rect 39304 44872 39356 44878
rect 39304 44814 39356 44820
rect 39672 44872 39724 44878
rect 39672 44814 39724 44820
rect 39120 44464 39172 44470
rect 39120 44406 39172 44412
rect 38936 43988 38988 43994
rect 38936 43930 38988 43936
rect 39132 43926 39160 44406
rect 39316 44402 39344 44814
rect 39304 44396 39356 44402
rect 39304 44338 39356 44344
rect 39684 44198 39712 44814
rect 39672 44192 39724 44198
rect 39672 44134 39724 44140
rect 39028 43920 39080 43926
rect 39026 43888 39028 43897
rect 39120 43920 39172 43926
rect 39080 43888 39082 43897
rect 39120 43862 39172 43868
rect 39026 43823 39082 43832
rect 38804 43744 38884 43772
rect 38936 43784 38988 43790
rect 38752 43726 38804 43732
rect 38936 43726 38988 43732
rect 38568 42696 38620 42702
rect 38568 42638 38620 42644
rect 38384 41812 38436 41818
rect 38384 41754 38436 41760
rect 38476 41132 38528 41138
rect 38476 41074 38528 41080
rect 38488 40186 38516 41074
rect 38580 40934 38608 42638
rect 38660 42628 38712 42634
rect 38660 42570 38712 42576
rect 38672 41478 38700 42570
rect 38948 42362 38976 43726
rect 39684 42634 39712 44134
rect 39776 43926 39804 45426
rect 40144 45404 40172 46514
rect 40500 45824 40552 45830
rect 40500 45766 40552 45772
rect 40512 45490 40540 45766
rect 40500 45484 40552 45490
rect 40500 45426 40552 45432
rect 40144 45376 40264 45404
rect 40132 44940 40184 44946
rect 40132 44882 40184 44888
rect 39856 44872 39908 44878
rect 39856 44814 39908 44820
rect 39868 44538 39896 44814
rect 39856 44532 39908 44538
rect 39856 44474 39908 44480
rect 39764 43920 39816 43926
rect 39764 43862 39816 43868
rect 39776 43790 39804 43862
rect 39764 43784 39816 43790
rect 39764 43726 39816 43732
rect 40040 43784 40092 43790
rect 40040 43726 40092 43732
rect 40052 42906 40080 43726
rect 40040 42900 40092 42906
rect 40040 42842 40092 42848
rect 39672 42628 39724 42634
rect 39672 42570 39724 42576
rect 38936 42356 38988 42362
rect 38936 42298 38988 42304
rect 39304 42288 39356 42294
rect 39304 42230 39356 42236
rect 39120 42220 39172 42226
rect 39120 42162 39172 42168
rect 38660 41472 38712 41478
rect 38660 41414 38712 41420
rect 39132 41274 39160 42162
rect 39316 41614 39344 42230
rect 39684 42022 39712 42570
rect 39672 42016 39724 42022
rect 39672 41958 39724 41964
rect 39304 41608 39356 41614
rect 39304 41550 39356 41556
rect 39948 41540 40000 41546
rect 39948 41482 40000 41488
rect 39960 41274 39988 41482
rect 39120 41268 39172 41274
rect 39120 41210 39172 41216
rect 39948 41268 40000 41274
rect 39948 41210 40000 41216
rect 38568 40928 38620 40934
rect 38568 40870 38620 40876
rect 38580 40526 38608 40870
rect 39960 40594 39988 41210
rect 39948 40588 40000 40594
rect 39948 40530 40000 40536
rect 38568 40520 38620 40526
rect 38568 40462 38620 40468
rect 39120 40520 39172 40526
rect 39120 40462 39172 40468
rect 39132 40390 39160 40462
rect 38752 40384 38804 40390
rect 38752 40326 38804 40332
rect 39120 40384 39172 40390
rect 39120 40326 39172 40332
rect 39488 40384 39540 40390
rect 39488 40326 39540 40332
rect 38476 40180 38528 40186
rect 38476 40122 38528 40128
rect 38384 40044 38436 40050
rect 38384 39986 38436 39992
rect 38396 38962 38424 39986
rect 38660 39500 38712 39506
rect 38660 39442 38712 39448
rect 38568 39296 38620 39302
rect 38568 39238 38620 39244
rect 38476 39092 38528 39098
rect 38476 39034 38528 39040
rect 38384 38956 38436 38962
rect 38384 38898 38436 38904
rect 38396 37777 38424 38898
rect 38488 38282 38516 39034
rect 38580 38962 38608 39238
rect 38568 38956 38620 38962
rect 38568 38898 38620 38904
rect 38672 38554 38700 39442
rect 38660 38548 38712 38554
rect 38660 38490 38712 38496
rect 38764 38418 38792 40326
rect 39500 40118 39528 40326
rect 39488 40112 39540 40118
rect 39488 40054 39540 40060
rect 39488 39976 39540 39982
rect 39856 39976 39908 39982
rect 39488 39918 39540 39924
rect 39684 39936 39856 39964
rect 39304 39432 39356 39438
rect 39304 39374 39356 39380
rect 39028 38820 39080 38826
rect 39028 38762 39080 38768
rect 38752 38412 38804 38418
rect 38752 38354 38804 38360
rect 38476 38276 38528 38282
rect 38476 38218 38528 38224
rect 38382 37768 38438 37777
rect 38382 37703 38438 37712
rect 38764 37398 38792 38354
rect 39040 38282 39068 38762
rect 39028 38276 39080 38282
rect 39028 38218 39080 38224
rect 38936 38208 38988 38214
rect 38936 38150 38988 38156
rect 38752 37392 38804 37398
rect 38752 37334 38804 37340
rect 38384 37120 38436 37126
rect 38384 37062 38436 37068
rect 38396 34678 38424 37062
rect 38764 35766 38792 37334
rect 38752 35760 38804 35766
rect 38752 35702 38804 35708
rect 38752 35488 38804 35494
rect 38752 35430 38804 35436
rect 38660 35080 38712 35086
rect 38660 35022 38712 35028
rect 38672 34746 38700 35022
rect 38660 34740 38712 34746
rect 38660 34682 38712 34688
rect 38384 34672 38436 34678
rect 38384 34614 38436 34620
rect 38672 34066 38700 34682
rect 38660 34060 38712 34066
rect 38660 34002 38712 34008
rect 38764 33998 38792 35430
rect 38752 33992 38804 33998
rect 38752 33934 38804 33940
rect 38752 32768 38804 32774
rect 38752 32710 38804 32716
rect 38660 32224 38712 32230
rect 38660 32166 38712 32172
rect 38304 31726 38424 31754
rect 38292 28960 38344 28966
rect 38292 28902 38344 28908
rect 38108 28416 38160 28422
rect 38108 28358 38160 28364
rect 37924 28076 37976 28082
rect 37924 28018 37976 28024
rect 37188 27940 37240 27946
rect 37188 27882 37240 27888
rect 37660 27934 37872 27962
rect 37200 27674 37228 27882
rect 37188 27668 37240 27674
rect 37188 27610 37240 27616
rect 37660 27470 37688 27934
rect 37844 27878 37872 27934
rect 37740 27872 37792 27878
rect 37740 27814 37792 27820
rect 37832 27872 37884 27878
rect 37832 27814 37884 27820
rect 37096 27464 37148 27470
rect 37096 27406 37148 27412
rect 37372 27464 37424 27470
rect 37372 27406 37424 27412
rect 37648 27464 37700 27470
rect 37648 27406 37700 27412
rect 37752 27452 37780 27814
rect 37936 27656 37964 28018
rect 38016 27668 38068 27674
rect 37936 27628 38016 27656
rect 38016 27610 38068 27616
rect 38120 27656 38148 28358
rect 38304 28218 38332 28902
rect 38292 28212 38344 28218
rect 38292 28154 38344 28160
rect 38200 27668 38252 27674
rect 38120 27628 38200 27656
rect 38016 27532 38068 27538
rect 38016 27474 38068 27480
rect 37832 27464 37884 27470
rect 37752 27424 37832 27452
rect 36820 27056 36872 27062
rect 36820 26998 36872 27004
rect 36728 26988 36780 26994
rect 36728 26930 36780 26936
rect 36544 26852 36596 26858
rect 36544 26794 36596 26800
rect 37108 26518 37136 27406
rect 37096 26512 37148 26518
rect 37096 26454 37148 26460
rect 37108 25362 37136 26454
rect 37280 26240 37332 26246
rect 37280 26182 37332 26188
rect 37292 25906 37320 26182
rect 37384 26042 37412 27406
rect 37752 27130 37780 27424
rect 37832 27406 37884 27412
rect 37740 27124 37792 27130
rect 37740 27066 37792 27072
rect 37832 26988 37884 26994
rect 37832 26930 37884 26936
rect 37648 26920 37700 26926
rect 37648 26862 37700 26868
rect 37372 26036 37424 26042
rect 37372 25978 37424 25984
rect 37280 25900 37332 25906
rect 37280 25842 37332 25848
rect 37096 25356 37148 25362
rect 37096 25298 37148 25304
rect 37280 25288 37332 25294
rect 37384 25276 37412 25978
rect 37660 25906 37688 26862
rect 37844 26382 37872 26930
rect 37832 26376 37884 26382
rect 37752 26336 37832 26364
rect 37556 25900 37608 25906
rect 37556 25842 37608 25848
rect 37648 25900 37700 25906
rect 37648 25842 37700 25848
rect 37332 25248 37412 25276
rect 37568 25786 37596 25842
rect 37752 25786 37780 26336
rect 37832 26318 37884 26324
rect 38028 25906 38056 27474
rect 38120 26246 38148 27628
rect 38200 27610 38252 27616
rect 38304 27402 38332 28154
rect 38396 28082 38424 31726
rect 38672 31346 38700 32166
rect 38660 31340 38712 31346
rect 38660 31282 38712 31288
rect 38764 31090 38792 32710
rect 38844 31952 38896 31958
rect 38844 31894 38896 31900
rect 38856 31142 38884 31894
rect 38580 31062 38792 31090
rect 38844 31136 38896 31142
rect 38844 31078 38896 31084
rect 38580 30682 38608 31062
rect 38948 30954 38976 38150
rect 39316 37466 39344 39374
rect 39396 39024 39448 39030
rect 39394 38992 39396 39001
rect 39448 38992 39450 39001
rect 39394 38927 39450 38936
rect 39500 38894 39528 39918
rect 39580 39636 39632 39642
rect 39580 39578 39632 39584
rect 39488 38888 39540 38894
rect 39394 38856 39450 38865
rect 39488 38830 39540 38836
rect 39394 38791 39396 38800
rect 39448 38791 39450 38800
rect 39396 38762 39448 38768
rect 39500 37942 39528 38830
rect 39592 38332 39620 39578
rect 39684 38826 39712 39936
rect 39856 39918 39908 39924
rect 40144 39846 40172 44882
rect 40236 40662 40264 45376
rect 40500 45348 40552 45354
rect 40500 45290 40552 45296
rect 40316 43852 40368 43858
rect 40316 43794 40368 43800
rect 40328 43625 40356 43794
rect 40314 43616 40370 43625
rect 40314 43551 40370 43560
rect 40224 40656 40276 40662
rect 40224 40598 40276 40604
rect 40408 40384 40460 40390
rect 40408 40326 40460 40332
rect 40316 40112 40368 40118
rect 40316 40054 40368 40060
rect 40132 39840 40184 39846
rect 40132 39782 40184 39788
rect 40132 39636 40184 39642
rect 40132 39578 40184 39584
rect 40040 39432 40092 39438
rect 40040 39374 40092 39380
rect 39948 39364 40000 39370
rect 39948 39306 40000 39312
rect 39960 38944 39988 39306
rect 40052 38962 40080 39374
rect 39868 38916 39988 38944
rect 40040 38956 40092 38962
rect 39672 38820 39724 38826
rect 39672 38762 39724 38768
rect 39684 38486 39712 38762
rect 39672 38480 39724 38486
rect 39672 38422 39724 38428
rect 39868 38350 39896 38916
rect 40040 38898 40092 38904
rect 40144 38826 40172 39578
rect 40224 39432 40276 39438
rect 40224 39374 40276 39380
rect 40236 39098 40264 39374
rect 40224 39092 40276 39098
rect 40224 39034 40276 39040
rect 40132 38820 40184 38826
rect 40132 38762 40184 38768
rect 40040 38412 40092 38418
rect 40040 38354 40092 38360
rect 39856 38344 39908 38350
rect 39592 38304 39712 38332
rect 39578 38040 39634 38049
rect 39578 37975 39580 37984
rect 39632 37975 39634 37984
rect 39580 37946 39632 37952
rect 39488 37936 39540 37942
rect 39488 37878 39540 37884
rect 39304 37460 39356 37466
rect 39304 37402 39356 37408
rect 39120 34944 39172 34950
rect 39120 34886 39172 34892
rect 39132 34202 39160 34886
rect 39120 34196 39172 34202
rect 39120 34138 39172 34144
rect 39120 33992 39172 33998
rect 39120 33934 39172 33940
rect 39132 33318 39160 33934
rect 39304 33856 39356 33862
rect 39304 33798 39356 33804
rect 39120 33312 39172 33318
rect 39120 33254 39172 33260
rect 39212 31476 39264 31482
rect 39212 31418 39264 31424
rect 39120 31204 39172 31210
rect 39120 31146 39172 31152
rect 39028 31136 39080 31142
rect 39028 31078 39080 31084
rect 38764 30926 38976 30954
rect 39040 30938 39068 31078
rect 39028 30932 39080 30938
rect 38580 30654 38700 30682
rect 38672 30394 38700 30654
rect 38660 30388 38712 30394
rect 38660 30330 38712 30336
rect 38764 30274 38792 30926
rect 39028 30874 39080 30880
rect 38936 30796 38988 30802
rect 38936 30738 38988 30744
rect 38844 30388 38896 30394
rect 38844 30330 38896 30336
rect 38672 30258 38792 30274
rect 38660 30252 38792 30258
rect 38712 30246 38792 30252
rect 38660 30194 38712 30200
rect 38568 30184 38620 30190
rect 38568 30126 38620 30132
rect 38476 29708 38528 29714
rect 38476 29650 38528 29656
rect 38488 29170 38516 29650
rect 38580 29322 38608 30126
rect 38672 29850 38700 30194
rect 38660 29844 38712 29850
rect 38660 29786 38712 29792
rect 38752 29844 38804 29850
rect 38752 29786 38804 29792
rect 38764 29646 38792 29786
rect 38752 29640 38804 29646
rect 38752 29582 38804 29588
rect 38580 29294 38700 29322
rect 38476 29164 38528 29170
rect 38476 29106 38528 29112
rect 38672 29034 38700 29294
rect 38856 29170 38884 30330
rect 38844 29164 38896 29170
rect 38844 29106 38896 29112
rect 38660 29028 38712 29034
rect 38660 28970 38712 28976
rect 38384 28076 38436 28082
rect 38384 28018 38436 28024
rect 38292 27396 38344 27402
rect 38292 27338 38344 27344
rect 38396 26994 38424 28018
rect 38856 27062 38884 29106
rect 38948 28558 38976 30738
rect 39132 30734 39160 31146
rect 39120 30728 39172 30734
rect 39120 30670 39172 30676
rect 39224 30546 39252 31418
rect 39316 30734 39344 33798
rect 39684 31482 39712 38304
rect 39856 38286 39908 38292
rect 39948 38344 40000 38350
rect 39948 38286 40000 38292
rect 39960 38010 39988 38286
rect 39948 38004 40000 38010
rect 39948 37946 40000 37952
rect 39764 37936 39816 37942
rect 39764 37878 39816 37884
rect 39672 31476 39724 31482
rect 39672 31418 39724 31424
rect 39396 31340 39448 31346
rect 39396 31282 39448 31288
rect 39408 30870 39436 31282
rect 39488 31136 39540 31142
rect 39488 31078 39540 31084
rect 39396 30864 39448 30870
rect 39396 30806 39448 30812
rect 39304 30728 39356 30734
rect 39304 30670 39356 30676
rect 39040 30518 39252 30546
rect 38936 28552 38988 28558
rect 38936 28494 38988 28500
rect 39040 27946 39068 30518
rect 39212 29504 39264 29510
rect 39212 29446 39264 29452
rect 39304 29504 39356 29510
rect 39304 29446 39356 29452
rect 39224 28218 39252 29446
rect 39212 28212 39264 28218
rect 39212 28154 39264 28160
rect 39212 28076 39264 28082
rect 39316 28064 39344 29446
rect 39264 28036 39344 28064
rect 39212 28018 39264 28024
rect 39028 27940 39080 27946
rect 39028 27882 39080 27888
rect 38844 27056 38896 27062
rect 38896 27016 38976 27044
rect 38844 26998 38896 27004
rect 38384 26988 38436 26994
rect 38384 26930 38436 26936
rect 38752 26784 38804 26790
rect 38752 26726 38804 26732
rect 38764 26450 38792 26726
rect 38752 26444 38804 26450
rect 38752 26386 38804 26392
rect 38660 26308 38712 26314
rect 38660 26250 38712 26256
rect 38108 26240 38160 26246
rect 38108 26182 38160 26188
rect 38016 25900 38068 25906
rect 38016 25842 38068 25848
rect 37568 25758 37780 25786
rect 37280 25230 37332 25236
rect 37568 24818 37596 25758
rect 38028 25294 38056 25842
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 37832 25152 37884 25158
rect 37832 25094 37884 25100
rect 37844 24886 37872 25094
rect 37832 24880 37884 24886
rect 37832 24822 37884 24828
rect 38120 24818 38148 26182
rect 38292 25696 38344 25702
rect 38292 25638 38344 25644
rect 38304 25294 38332 25638
rect 38292 25288 38344 25294
rect 38292 25230 38344 25236
rect 38672 24954 38700 26250
rect 38764 25838 38792 26386
rect 38844 26308 38896 26314
rect 38844 26250 38896 26256
rect 38856 25838 38884 26250
rect 38948 25906 38976 27016
rect 39224 26518 39252 28018
rect 39500 27334 39528 31078
rect 39776 29850 39804 37878
rect 39948 30728 40000 30734
rect 39948 30670 40000 30676
rect 39960 30258 39988 30670
rect 39948 30252 40000 30258
rect 39948 30194 40000 30200
rect 39764 29844 39816 29850
rect 39764 29786 39816 29792
rect 40052 29782 40080 38354
rect 40328 38214 40356 40054
rect 40420 39506 40448 40326
rect 40408 39500 40460 39506
rect 40408 39442 40460 39448
rect 40316 38208 40368 38214
rect 40316 38150 40368 38156
rect 40328 37874 40356 38150
rect 40420 37874 40448 39442
rect 40512 39098 40540 45290
rect 40592 44804 40644 44810
rect 40592 44746 40644 44752
rect 40604 44470 40632 44746
rect 40592 44464 40644 44470
rect 40592 44406 40644 44412
rect 40696 44033 40724 48486
rect 40960 48272 41012 48278
rect 40960 48214 41012 48220
rect 40868 48068 40920 48074
rect 40868 48010 40920 48016
rect 40880 47462 40908 48010
rect 40868 47456 40920 47462
rect 40868 47398 40920 47404
rect 40972 47258 41000 48214
rect 41052 48204 41104 48210
rect 41052 48146 41104 48152
rect 40960 47252 41012 47258
rect 40960 47194 41012 47200
rect 40866 47016 40922 47025
rect 40866 46951 40922 46960
rect 40880 46578 40908 46951
rect 41064 46714 41092 48146
rect 41156 48142 41184 48622
rect 41144 48136 41196 48142
rect 41144 48078 41196 48084
rect 41156 47666 41184 48078
rect 41144 47660 41196 47666
rect 41144 47602 41196 47608
rect 41420 47660 41472 47666
rect 41420 47602 41472 47608
rect 41328 47252 41380 47258
rect 41328 47194 41380 47200
rect 41340 47122 41368 47194
rect 41328 47116 41380 47122
rect 41328 47058 41380 47064
rect 41432 47054 41460 47602
rect 41420 47048 41472 47054
rect 41420 46990 41472 46996
rect 41052 46708 41104 46714
rect 41052 46650 41104 46656
rect 40868 46572 40920 46578
rect 40868 46514 40920 46520
rect 40776 45892 40828 45898
rect 40776 45834 40828 45840
rect 40788 45354 40816 45834
rect 40776 45348 40828 45354
rect 40776 45290 40828 45296
rect 40682 44024 40738 44033
rect 40682 43959 40738 43968
rect 40696 43790 40724 43959
rect 40684 43784 40736 43790
rect 40684 43726 40736 43732
rect 40684 41132 40736 41138
rect 40684 41074 40736 41080
rect 40592 40384 40644 40390
rect 40592 40326 40644 40332
rect 40604 40118 40632 40326
rect 40696 40186 40724 41074
rect 40788 40730 40816 45290
rect 40880 44538 40908 46514
rect 41064 46510 41092 46650
rect 41052 46504 41104 46510
rect 41052 46446 41104 46452
rect 41236 46096 41288 46102
rect 41236 46038 41288 46044
rect 41248 45490 41276 46038
rect 41236 45484 41288 45490
rect 41236 45426 41288 45432
rect 40960 45416 41012 45422
rect 40960 45358 41012 45364
rect 40972 45082 41000 45358
rect 40960 45076 41012 45082
rect 40960 45018 41012 45024
rect 41052 44872 41104 44878
rect 41052 44814 41104 44820
rect 40958 44704 41014 44713
rect 40958 44639 41014 44648
rect 40868 44532 40920 44538
rect 40868 44474 40920 44480
rect 40972 43654 41000 44639
rect 41064 44305 41092 44814
rect 41144 44396 41196 44402
rect 41144 44338 41196 44344
rect 41050 44296 41106 44305
rect 41050 44231 41106 44240
rect 41064 43722 41092 44231
rect 41156 43790 41184 44338
rect 41248 44266 41276 45426
rect 41328 45076 41380 45082
rect 41328 45018 41380 45024
rect 41340 44402 41368 45018
rect 41328 44396 41380 44402
rect 41328 44338 41380 44344
rect 41236 44260 41288 44266
rect 41236 44202 41288 44208
rect 41144 43784 41196 43790
rect 41144 43726 41196 43732
rect 41052 43716 41104 43722
rect 41052 43658 41104 43664
rect 40960 43648 41012 43654
rect 40960 43590 41012 43596
rect 40960 43104 41012 43110
rect 40960 43046 41012 43052
rect 40868 41064 40920 41070
rect 40868 41006 40920 41012
rect 40776 40724 40828 40730
rect 40776 40666 40828 40672
rect 40880 40594 40908 41006
rect 40868 40588 40920 40594
rect 40868 40530 40920 40536
rect 40684 40180 40736 40186
rect 40684 40122 40736 40128
rect 40592 40112 40644 40118
rect 40592 40054 40644 40060
rect 40880 39370 40908 40530
rect 40972 39642 41000 43046
rect 41156 42566 41184 43726
rect 41328 43648 41380 43654
rect 41328 43590 41380 43596
rect 41340 43450 41368 43590
rect 41328 43444 41380 43450
rect 41328 43386 41380 43392
rect 41236 43308 41288 43314
rect 41236 43250 41288 43256
rect 41248 42906 41276 43250
rect 41236 42900 41288 42906
rect 41236 42842 41288 42848
rect 41432 42702 41460 46990
rect 41524 46918 41552 49710
rect 48976 49298 49004 59200
rect 50264 57882 50292 59200
rect 50172 57854 50292 57882
rect 49700 56840 49752 56846
rect 49700 56782 49752 56788
rect 49712 56438 49740 56782
rect 49700 56432 49752 56438
rect 49700 56374 49752 56380
rect 50172 56234 50200 57854
rect 50294 57692 50602 57712
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57616 50602 57636
rect 55496 56840 55548 56846
rect 55496 56782 55548 56788
rect 50294 56604 50602 56624
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56528 50602 56548
rect 55508 56370 55536 56782
rect 55496 56364 55548 56370
rect 55496 56306 55548 56312
rect 50252 56296 50304 56302
rect 50252 56238 50304 56244
rect 50160 56228 50212 56234
rect 50160 56170 50212 56176
rect 50264 55962 50292 56238
rect 50252 55956 50304 55962
rect 50252 55898 50304 55904
rect 55404 55956 55456 55962
rect 55404 55898 55456 55904
rect 52920 55752 52972 55758
rect 52920 55694 52972 55700
rect 55312 55752 55364 55758
rect 55312 55694 55364 55700
rect 50294 55516 50602 55536
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55440 50602 55460
rect 52932 54534 52960 55694
rect 54668 55684 54720 55690
rect 54668 55626 54720 55632
rect 54680 55418 54708 55626
rect 54668 55412 54720 55418
rect 54668 55354 54720 55360
rect 55324 55350 55352 55694
rect 55312 55344 55364 55350
rect 55312 55286 55364 55292
rect 55416 55282 55444 55898
rect 56060 55826 56088 59200
rect 56506 58576 56562 58585
rect 56506 58511 56562 58520
rect 56324 57248 56376 57254
rect 56324 57190 56376 57196
rect 56336 56914 56364 57190
rect 56324 56908 56376 56914
rect 56324 56850 56376 56856
rect 56232 56160 56284 56166
rect 56232 56102 56284 56108
rect 56244 55894 56272 56102
rect 56232 55888 56284 55894
rect 56232 55830 56284 55836
rect 56520 55826 56548 58511
rect 56600 57248 56652 57254
rect 56600 57190 56652 57196
rect 56048 55820 56100 55826
rect 56048 55762 56100 55768
rect 56508 55820 56560 55826
rect 56508 55762 56560 55768
rect 55680 55752 55732 55758
rect 55680 55694 55732 55700
rect 55404 55276 55456 55282
rect 55404 55218 55456 55224
rect 52920 54528 52972 54534
rect 52920 54470 52972 54476
rect 50294 54428 50602 54448
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54352 50602 54372
rect 50294 53340 50602 53360
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53264 50602 53284
rect 50294 52252 50602 52272
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52176 50602 52196
rect 50294 51164 50602 51184
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51088 50602 51108
rect 50294 50076 50602 50096
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50000 50602 50020
rect 48964 49292 49016 49298
rect 48964 49234 49016 49240
rect 41788 49224 41840 49230
rect 41788 49166 41840 49172
rect 42708 49224 42760 49230
rect 42708 49166 42760 49172
rect 47768 49224 47820 49230
rect 47768 49166 47820 49172
rect 41800 48822 41828 49166
rect 41972 49156 42024 49162
rect 41972 49098 42024 49104
rect 41788 48816 41840 48822
rect 41788 48758 41840 48764
rect 41800 48210 41828 48758
rect 41880 48748 41932 48754
rect 41880 48690 41932 48696
rect 41892 48618 41920 48690
rect 41880 48612 41932 48618
rect 41880 48554 41932 48560
rect 41892 48346 41920 48554
rect 41880 48340 41932 48346
rect 41880 48282 41932 48288
rect 41788 48204 41840 48210
rect 41788 48146 41840 48152
rect 41984 48142 42012 49098
rect 42720 48686 42748 49166
rect 43536 49156 43588 49162
rect 43536 49098 43588 49104
rect 42892 49088 42944 49094
rect 42892 49030 42944 49036
rect 42524 48680 42576 48686
rect 42524 48622 42576 48628
rect 42708 48680 42760 48686
rect 42708 48622 42760 48628
rect 41972 48136 42024 48142
rect 41972 48078 42024 48084
rect 41696 47456 41748 47462
rect 41696 47398 41748 47404
rect 41512 46912 41564 46918
rect 41512 46854 41564 46860
rect 41524 46617 41552 46854
rect 41510 46608 41566 46617
rect 41510 46543 41566 46552
rect 41708 45966 41736 47398
rect 41970 47016 42026 47025
rect 41970 46951 41972 46960
rect 42024 46951 42026 46960
rect 42432 46980 42484 46986
rect 41972 46922 42024 46928
rect 42432 46922 42484 46928
rect 41696 45960 41748 45966
rect 41696 45902 41748 45908
rect 41696 45824 41748 45830
rect 41696 45766 41748 45772
rect 41604 45416 41656 45422
rect 41604 45358 41656 45364
rect 41708 45404 41736 45766
rect 41880 45416 41932 45422
rect 41708 45376 41880 45404
rect 41616 45014 41644 45358
rect 41604 45008 41656 45014
rect 41604 44950 41656 44956
rect 41708 44282 41736 45376
rect 41880 45358 41932 45364
rect 41788 44532 41840 44538
rect 41788 44474 41840 44480
rect 41524 44254 41736 44282
rect 41420 42696 41472 42702
rect 41420 42638 41472 42644
rect 41144 42560 41196 42566
rect 41144 42502 41196 42508
rect 41156 42226 41184 42502
rect 41144 42220 41196 42226
rect 41144 42162 41196 42168
rect 40960 39636 41012 39642
rect 40960 39578 41012 39584
rect 40592 39364 40644 39370
rect 40592 39306 40644 39312
rect 40868 39364 40920 39370
rect 40868 39306 40920 39312
rect 40500 39092 40552 39098
rect 40500 39034 40552 39040
rect 40604 38962 40632 39306
rect 40592 38956 40644 38962
rect 40592 38898 40644 38904
rect 40590 38856 40646 38865
rect 40590 38791 40646 38800
rect 40604 38758 40632 38791
rect 40592 38752 40644 38758
rect 40592 38694 40644 38700
rect 40684 38344 40736 38350
rect 40684 38286 40736 38292
rect 40696 37942 40724 38286
rect 40684 37936 40736 37942
rect 40684 37878 40736 37884
rect 40132 37868 40184 37874
rect 40132 37810 40184 37816
rect 40316 37868 40368 37874
rect 40316 37810 40368 37816
rect 40408 37868 40460 37874
rect 40408 37810 40460 37816
rect 40144 34202 40172 37810
rect 40328 36378 40356 37810
rect 40420 37262 40448 37810
rect 40682 37768 40738 37777
rect 40682 37703 40738 37712
rect 40592 37460 40644 37466
rect 40592 37402 40644 37408
rect 40604 37262 40632 37402
rect 40408 37256 40460 37262
rect 40592 37256 40644 37262
rect 40408 37198 40460 37204
rect 40512 37216 40592 37244
rect 40512 37108 40540 37216
rect 40592 37198 40644 37204
rect 40420 37080 40540 37108
rect 40592 37120 40644 37126
rect 40420 36854 40448 37080
rect 40592 37062 40644 37068
rect 40604 36854 40632 37062
rect 40408 36848 40460 36854
rect 40408 36790 40460 36796
rect 40592 36848 40644 36854
rect 40592 36790 40644 36796
rect 40500 36780 40552 36786
rect 40500 36722 40552 36728
rect 40316 36372 40368 36378
rect 40316 36314 40368 36320
rect 40408 35692 40460 35698
rect 40408 35634 40460 35640
rect 40420 34746 40448 35634
rect 40408 34740 40460 34746
rect 40408 34682 40460 34688
rect 40316 34672 40368 34678
rect 40316 34614 40368 34620
rect 40132 34196 40184 34202
rect 40132 34138 40184 34144
rect 40328 31482 40356 34614
rect 40408 34604 40460 34610
rect 40408 34546 40460 34552
rect 40420 34513 40448 34546
rect 40512 34542 40540 36722
rect 40500 34536 40552 34542
rect 40406 34504 40462 34513
rect 40500 34478 40552 34484
rect 40406 34439 40462 34448
rect 40316 31476 40368 31482
rect 40316 31418 40368 31424
rect 40224 30592 40276 30598
rect 40224 30534 40276 30540
rect 40236 29782 40264 30534
rect 40328 30394 40356 31418
rect 40408 30660 40460 30666
rect 40408 30602 40460 30608
rect 40316 30388 40368 30394
rect 40316 30330 40368 30336
rect 40316 30048 40368 30054
rect 40316 29990 40368 29996
rect 40040 29776 40092 29782
rect 40040 29718 40092 29724
rect 40224 29776 40276 29782
rect 40224 29718 40276 29724
rect 40052 29628 40080 29718
rect 40132 29640 40184 29646
rect 40052 29600 40132 29628
rect 40132 29582 40184 29588
rect 39580 29572 39632 29578
rect 39580 29514 39632 29520
rect 40224 29572 40276 29578
rect 40224 29514 40276 29520
rect 39592 29238 39620 29514
rect 39580 29232 39632 29238
rect 39580 29174 39632 29180
rect 40236 28490 40264 29514
rect 40224 28484 40276 28490
rect 40224 28426 40276 28432
rect 39488 27328 39540 27334
rect 39488 27270 39540 27276
rect 40224 26920 40276 26926
rect 40224 26862 40276 26868
rect 40040 26852 40092 26858
rect 40040 26794 40092 26800
rect 39212 26512 39264 26518
rect 39212 26454 39264 26460
rect 40052 26382 40080 26794
rect 40040 26376 40092 26382
rect 40040 26318 40092 26324
rect 39764 26240 39816 26246
rect 39764 26182 39816 26188
rect 39580 25968 39632 25974
rect 39578 25936 39580 25945
rect 39632 25936 39634 25945
rect 38936 25900 38988 25906
rect 38936 25842 38988 25848
rect 39488 25900 39540 25906
rect 39578 25871 39634 25880
rect 39776 25922 39804 26182
rect 39856 25934 39908 25940
rect 39776 25894 39856 25922
rect 39488 25842 39540 25848
rect 38752 25832 38804 25838
rect 38752 25774 38804 25780
rect 38844 25832 38896 25838
rect 38844 25774 38896 25780
rect 38764 25430 38792 25774
rect 38752 25424 38804 25430
rect 38752 25366 38804 25372
rect 38856 25294 38884 25774
rect 39120 25424 39172 25430
rect 39120 25366 39172 25372
rect 39132 25294 39160 25366
rect 39500 25362 39528 25842
rect 39488 25356 39540 25362
rect 39488 25298 39540 25304
rect 38844 25288 38896 25294
rect 38844 25230 38896 25236
rect 39120 25288 39172 25294
rect 39120 25230 39172 25236
rect 39776 25226 39804 25894
rect 39856 25876 39908 25882
rect 40040 25900 40092 25906
rect 40092 25860 40172 25888
rect 40040 25842 40092 25848
rect 40040 25492 40092 25498
rect 40040 25434 40092 25440
rect 39764 25220 39816 25226
rect 39764 25162 39816 25168
rect 39120 25152 39172 25158
rect 39120 25094 39172 25100
rect 38660 24948 38712 24954
rect 38660 24890 38712 24896
rect 38844 24948 38896 24954
rect 38844 24890 38896 24896
rect 37556 24812 37608 24818
rect 37556 24754 37608 24760
rect 38108 24812 38160 24818
rect 38108 24754 38160 24760
rect 38672 24682 38700 24890
rect 38856 24818 38884 24890
rect 39132 24818 39160 25094
rect 38844 24812 38896 24818
rect 38844 24754 38896 24760
rect 39120 24812 39172 24818
rect 39120 24754 39172 24760
rect 38660 24676 38712 24682
rect 38660 24618 38712 24624
rect 39304 24608 39356 24614
rect 39304 24550 39356 24556
rect 39316 24206 39344 24550
rect 39304 24200 39356 24206
rect 39304 24142 39356 24148
rect 40052 23254 40080 25434
rect 40144 25430 40172 25860
rect 40132 25424 40184 25430
rect 40132 25366 40184 25372
rect 40236 25158 40264 26862
rect 40328 26518 40356 29990
rect 40420 29782 40448 30602
rect 40512 30190 40540 34478
rect 40604 30598 40632 36790
rect 40696 34513 40724 37703
rect 40682 34504 40738 34513
rect 40682 34439 40738 34448
rect 40880 33862 40908 39306
rect 41156 37942 41184 42162
rect 41524 41414 41552 44254
rect 41696 43648 41748 43654
rect 41696 43590 41748 43596
rect 41604 42832 41656 42838
rect 41604 42774 41656 42780
rect 41616 42673 41644 42774
rect 41602 42664 41658 42673
rect 41602 42599 41658 42608
rect 41708 42158 41736 43590
rect 41800 43314 41828 44474
rect 41880 44396 41932 44402
rect 41880 44338 41932 44344
rect 41788 43308 41840 43314
rect 41788 43250 41840 43256
rect 41788 42832 41840 42838
rect 41788 42774 41840 42780
rect 41696 42152 41748 42158
rect 41696 42094 41748 42100
rect 41432 41386 41552 41414
rect 41432 41138 41460 41386
rect 41708 41274 41736 42094
rect 41696 41268 41748 41274
rect 41696 41210 41748 41216
rect 41800 41138 41828 42774
rect 41892 42226 41920 44338
rect 41984 44266 42012 46922
rect 42248 46572 42300 46578
rect 42248 46514 42300 46520
rect 42260 45898 42288 46514
rect 42248 45892 42300 45898
rect 42248 45834 42300 45840
rect 42156 45824 42208 45830
rect 42156 45766 42208 45772
rect 42064 45620 42116 45626
rect 42064 45562 42116 45568
rect 41972 44260 42024 44266
rect 41972 44202 42024 44208
rect 41984 43858 42012 44202
rect 41972 43852 42024 43858
rect 41972 43794 42024 43800
rect 42076 42786 42104 45562
rect 42168 43926 42196 45766
rect 42260 44810 42288 45834
rect 42444 45286 42472 46922
rect 42432 45280 42484 45286
rect 42432 45222 42484 45228
rect 42432 44872 42484 44878
rect 42432 44814 42484 44820
rect 42248 44804 42300 44810
rect 42248 44746 42300 44752
rect 42340 44736 42392 44742
rect 42444 44713 42472 44814
rect 42536 44742 42564 48622
rect 42904 48074 42932 49030
rect 42892 48068 42944 48074
rect 42892 48010 42944 48016
rect 42892 47048 42944 47054
rect 42892 46990 42944 46996
rect 42800 46980 42852 46986
rect 42800 46922 42852 46928
rect 42812 46578 42840 46922
rect 42904 46646 42932 46990
rect 43168 46912 43220 46918
rect 43168 46854 43220 46860
rect 42892 46640 42944 46646
rect 42892 46582 42944 46588
rect 42800 46572 42852 46578
rect 42800 46514 42852 46520
rect 42708 46368 42760 46374
rect 42708 46310 42760 46316
rect 42720 46170 42748 46310
rect 42708 46164 42760 46170
rect 42708 46106 42760 46112
rect 42720 45966 42748 46106
rect 42812 45966 42840 46514
rect 42904 46034 42932 46582
rect 43180 46102 43208 46854
rect 43352 46708 43404 46714
rect 43352 46650 43404 46656
rect 43168 46096 43220 46102
rect 43168 46038 43220 46044
rect 42892 46028 42944 46034
rect 42892 45970 42944 45976
rect 42708 45960 42760 45966
rect 42708 45902 42760 45908
rect 42800 45960 42852 45966
rect 42800 45902 42852 45908
rect 42984 45960 43036 45966
rect 42984 45902 43036 45908
rect 42812 45558 42840 45902
rect 42800 45552 42852 45558
rect 42800 45494 42852 45500
rect 42892 45484 42944 45490
rect 42996 45472 43024 45902
rect 43076 45824 43128 45830
rect 43076 45766 43128 45772
rect 42944 45444 43024 45472
rect 42892 45426 42944 45432
rect 43088 45422 43116 45766
rect 43180 45558 43208 46038
rect 43364 45898 43392 46650
rect 43352 45892 43404 45898
rect 43352 45834 43404 45840
rect 43168 45552 43220 45558
rect 43168 45494 43220 45500
rect 43076 45416 43128 45422
rect 43076 45358 43128 45364
rect 42892 44804 42944 44810
rect 42892 44746 42944 44752
rect 42984 44804 43036 44810
rect 42984 44746 43036 44752
rect 42524 44736 42576 44742
rect 42340 44678 42392 44684
rect 42430 44704 42486 44713
rect 42156 43920 42208 43926
rect 42156 43862 42208 43868
rect 42156 43240 42208 43246
rect 42154 43208 42156 43217
rect 42248 43240 42300 43246
rect 42208 43208 42210 43217
rect 42248 43182 42300 43188
rect 42154 43143 42210 43152
rect 42260 42906 42288 43182
rect 42248 42900 42300 42906
rect 42248 42842 42300 42848
rect 42076 42758 42288 42786
rect 42064 42696 42116 42702
rect 42064 42638 42116 42644
rect 42076 42362 42104 42638
rect 42064 42356 42116 42362
rect 42064 42298 42116 42304
rect 41880 42220 41932 42226
rect 41880 42162 41932 42168
rect 41420 41132 41472 41138
rect 41420 41074 41472 41080
rect 41604 41132 41656 41138
rect 41604 41074 41656 41080
rect 41788 41132 41840 41138
rect 41788 41074 41840 41080
rect 41432 39846 41460 41074
rect 41616 40526 41644 41074
rect 41696 40996 41748 41002
rect 41696 40938 41748 40944
rect 41708 40526 41736 40938
rect 41604 40520 41656 40526
rect 41604 40462 41656 40468
rect 41696 40520 41748 40526
rect 41696 40462 41748 40468
rect 41512 40384 41564 40390
rect 41512 40326 41564 40332
rect 41524 40050 41552 40326
rect 41512 40044 41564 40050
rect 41512 39986 41564 39992
rect 41420 39840 41472 39846
rect 41420 39782 41472 39788
rect 41326 38992 41382 39001
rect 41524 38962 41552 39986
rect 41616 39642 41644 40462
rect 41604 39636 41656 39642
rect 41604 39578 41656 39584
rect 41604 39024 41656 39030
rect 41604 38966 41656 38972
rect 41326 38927 41382 38936
rect 41512 38956 41564 38962
rect 41340 38554 41368 38927
rect 41512 38898 41564 38904
rect 41328 38548 41380 38554
rect 41328 38490 41380 38496
rect 41512 38344 41564 38350
rect 41512 38286 41564 38292
rect 41236 38208 41288 38214
rect 41236 38150 41288 38156
rect 41248 38010 41276 38150
rect 41236 38004 41288 38010
rect 41236 37946 41288 37952
rect 41144 37936 41196 37942
rect 41144 37878 41196 37884
rect 41052 37664 41104 37670
rect 41052 37606 41104 37612
rect 41064 37262 41092 37606
rect 41420 37392 41472 37398
rect 41420 37334 41472 37340
rect 41052 37256 41104 37262
rect 41052 37198 41104 37204
rect 41144 37256 41196 37262
rect 41144 37198 41196 37204
rect 40960 35488 41012 35494
rect 40960 35430 41012 35436
rect 40972 35154 41000 35430
rect 41064 35290 41092 37198
rect 41156 36854 41184 37198
rect 41432 36854 41460 37334
rect 41524 37126 41552 38286
rect 41616 38282 41644 38966
rect 41800 38593 41828 41074
rect 42260 40526 42288 42758
rect 42352 41546 42380 44678
rect 42524 44678 42576 44684
rect 42430 44639 42486 44648
rect 42444 43790 42472 44639
rect 42904 44402 42932 44746
rect 42996 44538 43024 44746
rect 42984 44532 43036 44538
rect 42984 44474 43036 44480
rect 42892 44396 42944 44402
rect 42892 44338 42944 44344
rect 42708 44260 42760 44266
rect 42708 44202 42760 44208
rect 42432 43784 42484 43790
rect 42432 43726 42484 43732
rect 42616 43648 42668 43654
rect 42616 43590 42668 43596
rect 42628 43450 42656 43590
rect 42616 43444 42668 43450
rect 42616 43386 42668 43392
rect 42524 43308 42576 43314
rect 42524 43250 42576 43256
rect 42432 42288 42484 42294
rect 42432 42230 42484 42236
rect 42444 42090 42472 42230
rect 42432 42084 42484 42090
rect 42432 42026 42484 42032
rect 42536 41750 42564 43250
rect 42720 42906 42748 44202
rect 42800 44192 42852 44198
rect 42800 44134 42852 44140
rect 42812 43722 42840 44134
rect 42982 43888 43038 43897
rect 42982 43823 43038 43832
rect 42996 43722 43024 43823
rect 42800 43716 42852 43722
rect 42800 43658 42852 43664
rect 42984 43716 43036 43722
rect 42984 43658 43036 43664
rect 42892 43648 42944 43654
rect 42892 43590 42944 43596
rect 42904 43450 42932 43590
rect 42982 43480 43038 43489
rect 42800 43444 42852 43450
rect 42800 43386 42852 43392
rect 42892 43444 42944 43450
rect 42982 43415 43038 43424
rect 42892 43386 42944 43392
rect 42708 42900 42760 42906
rect 42812 42888 42840 43386
rect 42892 43308 42944 43314
rect 42996 43296 43024 43415
rect 42944 43268 43024 43296
rect 42892 43250 42944 43256
rect 43088 43178 43116 45358
rect 43168 44804 43220 44810
rect 43168 44746 43220 44752
rect 43180 44402 43208 44746
rect 43168 44396 43220 44402
rect 43168 44338 43220 44344
rect 43260 44328 43312 44334
rect 43260 44270 43312 44276
rect 43168 43308 43220 43314
rect 43168 43250 43220 43256
rect 43076 43172 43128 43178
rect 43076 43114 43128 43120
rect 42812 42860 42932 42888
rect 42708 42842 42760 42848
rect 42800 42764 42852 42770
rect 42800 42706 42852 42712
rect 42812 42362 42840 42706
rect 42904 42566 42932 42860
rect 43088 42634 43116 43114
rect 43076 42628 43128 42634
rect 43076 42570 43128 42576
rect 42892 42560 42944 42566
rect 42892 42502 42944 42508
rect 42800 42356 42852 42362
rect 42800 42298 42852 42304
rect 42708 42016 42760 42022
rect 42708 41958 42760 41964
rect 42524 41744 42576 41750
rect 42524 41686 42576 41692
rect 42432 41608 42484 41614
rect 42432 41550 42484 41556
rect 42340 41540 42392 41546
rect 42340 41482 42392 41488
rect 42444 41070 42472 41550
rect 42616 41472 42668 41478
rect 42616 41414 42668 41420
rect 42432 41064 42484 41070
rect 42432 41006 42484 41012
rect 42156 40520 42208 40526
rect 42156 40462 42208 40468
rect 42248 40520 42300 40526
rect 42248 40462 42300 40468
rect 41880 39636 41932 39642
rect 41880 39578 41932 39584
rect 41786 38584 41842 38593
rect 41786 38519 41842 38528
rect 41696 38480 41748 38486
rect 41696 38422 41748 38428
rect 41604 38276 41656 38282
rect 41604 38218 41656 38224
rect 41708 37992 41736 38422
rect 41616 37964 41736 37992
rect 41616 37874 41644 37964
rect 41604 37868 41656 37874
rect 41604 37810 41656 37816
rect 41512 37120 41564 37126
rect 41512 37062 41564 37068
rect 41144 36848 41196 36854
rect 41144 36790 41196 36796
rect 41420 36848 41472 36854
rect 41420 36790 41472 36796
rect 41696 36032 41748 36038
rect 41696 35974 41748 35980
rect 41708 35630 41736 35974
rect 41512 35624 41564 35630
rect 41512 35566 41564 35572
rect 41696 35624 41748 35630
rect 41696 35566 41748 35572
rect 41328 35488 41380 35494
rect 41328 35430 41380 35436
rect 41052 35284 41104 35290
rect 41052 35226 41104 35232
rect 40960 35148 41012 35154
rect 40960 35090 41012 35096
rect 41052 35148 41104 35154
rect 41052 35090 41104 35096
rect 41064 34066 41092 35090
rect 41340 35086 41368 35430
rect 41328 35080 41380 35086
rect 41328 35022 41380 35028
rect 41340 34678 41368 35022
rect 41420 34944 41472 34950
rect 41420 34886 41472 34892
rect 41328 34672 41380 34678
rect 41328 34614 41380 34620
rect 41432 34610 41460 34886
rect 41524 34746 41552 35566
rect 41512 34740 41564 34746
rect 41512 34682 41564 34688
rect 41524 34610 41552 34682
rect 41420 34604 41472 34610
rect 41420 34546 41472 34552
rect 41512 34604 41564 34610
rect 41512 34546 41564 34552
rect 41052 34060 41104 34066
rect 41052 34002 41104 34008
rect 40684 33856 40736 33862
rect 40684 33798 40736 33804
rect 40868 33856 40920 33862
rect 40868 33798 40920 33804
rect 41236 33856 41288 33862
rect 41236 33798 41288 33804
rect 40696 32570 40724 33798
rect 41248 33454 41276 33798
rect 41328 33584 41380 33590
rect 41328 33526 41380 33532
rect 41236 33448 41288 33454
rect 41236 33390 41288 33396
rect 41340 33114 41368 33526
rect 41328 33108 41380 33114
rect 41328 33050 41380 33056
rect 41236 32836 41288 32842
rect 41236 32778 41288 32784
rect 40684 32564 40736 32570
rect 40684 32506 40736 32512
rect 41248 32434 41276 32778
rect 41236 32428 41288 32434
rect 41236 32370 41288 32376
rect 41432 32026 41460 34546
rect 41604 34060 41656 34066
rect 41604 34002 41656 34008
rect 41616 33658 41644 34002
rect 41604 33652 41656 33658
rect 41604 33594 41656 33600
rect 41512 32904 41564 32910
rect 41512 32846 41564 32852
rect 41604 32904 41656 32910
rect 41604 32846 41656 32852
rect 41524 32434 41552 32846
rect 41616 32774 41644 32846
rect 41604 32768 41656 32774
rect 41604 32710 41656 32716
rect 41616 32570 41644 32710
rect 41604 32564 41656 32570
rect 41604 32506 41656 32512
rect 41708 32502 41736 35566
rect 41892 35290 41920 39578
rect 42168 39030 42196 40462
rect 42260 40050 42288 40462
rect 42248 40044 42300 40050
rect 42248 39986 42300 39992
rect 42156 39024 42208 39030
rect 42156 38966 42208 38972
rect 42444 38418 42472 41006
rect 42432 38412 42484 38418
rect 42432 38354 42484 38360
rect 42064 37868 42116 37874
rect 42064 37810 42116 37816
rect 42432 37868 42484 37874
rect 42432 37810 42484 37816
rect 42076 37466 42104 37810
rect 42156 37800 42208 37806
rect 42156 37742 42208 37748
rect 42168 37466 42196 37742
rect 42064 37460 42116 37466
rect 42064 37402 42116 37408
rect 42156 37460 42208 37466
rect 42156 37402 42208 37408
rect 42168 37194 42196 37402
rect 42444 37262 42472 37810
rect 42432 37256 42484 37262
rect 42432 37198 42484 37204
rect 42156 37188 42208 37194
rect 42156 37130 42208 37136
rect 41880 35284 41932 35290
rect 41880 35226 41932 35232
rect 42522 35184 42578 35193
rect 42522 35119 42524 35128
rect 42576 35119 42578 35128
rect 42524 35090 42576 35096
rect 41972 34400 42024 34406
rect 41972 34342 42024 34348
rect 41984 34066 42012 34342
rect 41972 34060 42024 34066
rect 41972 34002 42024 34008
rect 41880 33992 41932 33998
rect 41880 33934 41932 33940
rect 41892 33522 41920 33934
rect 42524 33924 42576 33930
rect 42524 33866 42576 33872
rect 41880 33516 41932 33522
rect 41880 33458 41932 33464
rect 42432 33516 42484 33522
rect 42432 33458 42484 33464
rect 42444 32570 42472 33458
rect 42536 33046 42564 33866
rect 42524 33040 42576 33046
rect 42524 32982 42576 32988
rect 42628 32774 42656 41414
rect 42720 40730 42748 41958
rect 43180 41614 43208 43250
rect 43272 42226 43300 44270
rect 43260 42220 43312 42226
rect 43260 42162 43312 42168
rect 43272 41818 43300 42162
rect 43260 41812 43312 41818
rect 43260 41754 43312 41760
rect 43168 41608 43220 41614
rect 43168 41550 43220 41556
rect 42892 41540 42944 41546
rect 42892 41482 42944 41488
rect 42904 41138 42932 41482
rect 42892 41132 42944 41138
rect 42892 41074 42944 41080
rect 42708 40724 42760 40730
rect 42708 40666 42760 40672
rect 42720 40458 42748 40666
rect 42904 40526 42932 41074
rect 43180 40594 43208 41550
rect 43168 40588 43220 40594
rect 43168 40530 43220 40536
rect 42892 40520 42944 40526
rect 42892 40462 42944 40468
rect 42708 40452 42760 40458
rect 42708 40394 42760 40400
rect 42708 40044 42760 40050
rect 42708 39986 42760 39992
rect 42720 37398 42748 39986
rect 42798 37904 42854 37913
rect 42798 37839 42800 37848
rect 42852 37839 42854 37848
rect 42800 37810 42852 37816
rect 42708 37392 42760 37398
rect 42708 37334 42760 37340
rect 42720 36650 42748 37334
rect 42708 36644 42760 36650
rect 42708 36586 42760 36592
rect 43168 36168 43220 36174
rect 43168 36110 43220 36116
rect 43180 35834 43208 36110
rect 43168 35828 43220 35834
rect 43168 35770 43220 35776
rect 43364 35766 43392 45834
rect 43444 45620 43496 45626
rect 43444 45562 43496 45568
rect 43456 45082 43484 45562
rect 43444 45076 43496 45082
rect 43444 45018 43496 45024
rect 43444 44532 43496 44538
rect 43444 44474 43496 44480
rect 43456 42226 43484 44474
rect 43548 44334 43576 49098
rect 44456 49088 44508 49094
rect 44456 49030 44508 49036
rect 43996 48544 44048 48550
rect 43996 48486 44048 48492
rect 44008 48142 44036 48486
rect 44088 48204 44140 48210
rect 44088 48146 44140 48152
rect 44272 48204 44324 48210
rect 44272 48146 44324 48152
rect 43996 48136 44048 48142
rect 43996 48078 44048 48084
rect 43628 48000 43680 48006
rect 43628 47942 43680 47948
rect 43640 46578 43668 47942
rect 44100 47734 44128 48146
rect 44088 47728 44140 47734
rect 44088 47670 44140 47676
rect 43628 46572 43680 46578
rect 43628 46514 43680 46520
rect 43904 46572 43956 46578
rect 43904 46514 43956 46520
rect 43640 45966 43668 46514
rect 43916 46034 43944 46514
rect 43904 46028 43956 46034
rect 43904 45970 43956 45976
rect 43628 45960 43680 45966
rect 43628 45902 43680 45908
rect 43536 44328 43588 44334
rect 43536 44270 43588 44276
rect 43444 42220 43496 42226
rect 43444 42162 43496 42168
rect 43456 41274 43484 42162
rect 43444 41268 43496 41274
rect 43444 41210 43496 41216
rect 43548 38894 43576 44270
rect 43640 43489 43668 45902
rect 44100 44878 44128 47670
rect 44180 47660 44232 47666
rect 44180 47602 44232 47608
rect 44192 47530 44220 47602
rect 44284 47598 44312 48146
rect 44272 47592 44324 47598
rect 44272 47534 44324 47540
rect 44180 47524 44232 47530
rect 44180 47466 44232 47472
rect 44192 46986 44220 47466
rect 44180 46980 44232 46986
rect 44180 46922 44232 46928
rect 44180 46504 44232 46510
rect 44180 46446 44232 46452
rect 44192 45966 44220 46446
rect 44468 45966 44496 49030
rect 47780 48890 47808 49166
rect 48228 49156 48280 49162
rect 48228 49098 48280 49104
rect 48240 48890 48268 49098
rect 50294 48988 50602 49008
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48912 50602 48932
rect 47768 48884 47820 48890
rect 47768 48826 47820 48832
rect 48228 48884 48280 48890
rect 48228 48826 48280 48832
rect 44916 48748 44968 48754
rect 44916 48690 44968 48696
rect 45008 48748 45060 48754
rect 45008 48690 45060 48696
rect 45192 48748 45244 48754
rect 45192 48690 45244 48696
rect 48136 48748 48188 48754
rect 48136 48690 48188 48696
rect 44928 47802 44956 48690
rect 44916 47796 44968 47802
rect 44916 47738 44968 47744
rect 44916 47660 44968 47666
rect 44916 47602 44968 47608
rect 44928 47122 44956 47602
rect 44916 47116 44968 47122
rect 44916 47058 44968 47064
rect 44732 46912 44784 46918
rect 44732 46854 44784 46860
rect 44744 46646 44772 46854
rect 44732 46640 44784 46646
rect 44732 46582 44784 46588
rect 45020 46170 45048 48690
rect 45204 48226 45232 48690
rect 46020 48680 46072 48686
rect 46020 48622 46072 48628
rect 45284 48544 45336 48550
rect 45284 48486 45336 48492
rect 45296 48278 45324 48486
rect 46032 48346 46060 48622
rect 46020 48340 46072 48346
rect 46020 48282 46072 48288
rect 48148 48278 48176 48690
rect 45112 48198 45232 48226
rect 45284 48272 45336 48278
rect 45284 48214 45336 48220
rect 48136 48272 48188 48278
rect 48136 48214 48188 48220
rect 46572 48204 46624 48210
rect 45112 46714 45140 48198
rect 46572 48146 46624 48152
rect 45192 48136 45244 48142
rect 45376 48136 45428 48142
rect 45192 48078 45244 48084
rect 45296 48096 45376 48124
rect 45204 47802 45232 48078
rect 45192 47796 45244 47802
rect 45192 47738 45244 47744
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 46708 45152 46714
rect 45100 46650 45152 46656
rect 45204 46578 45232 46990
rect 45192 46572 45244 46578
rect 45192 46514 45244 46520
rect 45296 46510 45324 48096
rect 45376 48078 45428 48084
rect 46296 48136 46348 48142
rect 46296 48078 46348 48084
rect 45836 48068 45888 48074
rect 45836 48010 45888 48016
rect 45468 48000 45520 48006
rect 45468 47942 45520 47948
rect 45480 47666 45508 47942
rect 45376 47660 45428 47666
rect 45376 47602 45428 47608
rect 45468 47660 45520 47666
rect 45468 47602 45520 47608
rect 45652 47660 45704 47666
rect 45652 47602 45704 47608
rect 45388 47258 45416 47602
rect 45376 47252 45428 47258
rect 45376 47194 45428 47200
rect 45376 47048 45428 47054
rect 45374 47016 45376 47025
rect 45428 47016 45430 47025
rect 45374 46951 45430 46960
rect 45560 46572 45612 46578
rect 45560 46514 45612 46520
rect 45284 46504 45336 46510
rect 45284 46446 45336 46452
rect 45008 46164 45060 46170
rect 45008 46106 45060 46112
rect 45572 46102 45600 46514
rect 45560 46096 45612 46102
rect 45560 46038 45612 46044
rect 44180 45960 44232 45966
rect 44180 45902 44232 45908
rect 44456 45960 44508 45966
rect 44456 45902 44508 45908
rect 44916 45960 44968 45966
rect 44916 45902 44968 45908
rect 44548 45892 44600 45898
rect 44548 45834 44600 45840
rect 44088 44872 44140 44878
rect 44088 44814 44140 44820
rect 44180 44804 44232 44810
rect 44180 44746 44232 44752
rect 44192 44538 44220 44746
rect 44364 44736 44416 44742
rect 44364 44678 44416 44684
rect 44180 44532 44232 44538
rect 44180 44474 44232 44480
rect 44376 44470 44404 44678
rect 44364 44464 44416 44470
rect 44364 44406 44416 44412
rect 43904 44396 43956 44402
rect 43904 44338 43956 44344
rect 43720 44328 43772 44334
rect 43720 44270 43772 44276
rect 43732 43994 43760 44270
rect 43720 43988 43772 43994
rect 43720 43930 43772 43936
rect 43626 43480 43682 43489
rect 43626 43415 43682 43424
rect 43916 41414 43944 44338
rect 44180 43784 44232 43790
rect 44180 43726 44232 43732
rect 43996 43648 44048 43654
rect 43996 43590 44048 43596
rect 44008 43314 44036 43590
rect 43996 43308 44048 43314
rect 43996 43250 44048 43256
rect 44088 43308 44140 43314
rect 44088 43250 44140 43256
rect 44100 43217 44128 43250
rect 44086 43208 44142 43217
rect 44086 43143 44142 43152
rect 43916 41386 44036 41414
rect 43536 38888 43588 38894
rect 43536 38830 43588 38836
rect 43536 38276 43588 38282
rect 43536 38218 43588 38224
rect 43720 38276 43772 38282
rect 43720 38218 43772 38224
rect 43548 38010 43576 38218
rect 43536 38004 43588 38010
rect 43536 37946 43588 37952
rect 43536 37868 43588 37874
rect 43732 37856 43760 38218
rect 43588 37828 43760 37856
rect 43536 37810 43588 37816
rect 43444 37120 43496 37126
rect 43444 37062 43496 37068
rect 43456 36378 43484 37062
rect 43444 36372 43496 36378
rect 43444 36314 43496 36320
rect 43536 36032 43588 36038
rect 43536 35974 43588 35980
rect 43352 35760 43404 35766
rect 43352 35702 43404 35708
rect 43444 35760 43496 35766
rect 43444 35702 43496 35708
rect 42892 35488 42944 35494
rect 42892 35430 42944 35436
rect 42708 35284 42760 35290
rect 42708 35226 42760 35232
rect 42720 33538 42748 35226
rect 42904 35222 42932 35430
rect 42892 35216 42944 35222
rect 42892 35158 42944 35164
rect 42904 34678 42932 35158
rect 43364 35154 43392 35702
rect 43352 35148 43404 35154
rect 43352 35090 43404 35096
rect 43260 35012 43312 35018
rect 43260 34954 43312 34960
rect 42800 34672 42852 34678
rect 42798 34640 42800 34649
rect 42892 34672 42944 34678
rect 42852 34640 42854 34649
rect 42892 34614 42944 34620
rect 42798 34575 42854 34584
rect 42984 33992 43036 33998
rect 42984 33934 43036 33940
rect 42800 33856 42852 33862
rect 42800 33798 42852 33804
rect 42812 33658 42840 33798
rect 42996 33658 43024 33934
rect 42800 33652 42852 33658
rect 42800 33594 42852 33600
rect 42984 33652 43036 33658
rect 42984 33594 43036 33600
rect 42892 33584 42944 33590
rect 42720 33532 42892 33538
rect 42720 33526 42944 33532
rect 42720 33510 42932 33526
rect 42708 33448 42760 33454
rect 42708 33390 42760 33396
rect 42720 33114 42748 33390
rect 42708 33108 42760 33114
rect 42708 33050 42760 33056
rect 42616 32768 42668 32774
rect 42616 32710 42668 32716
rect 42432 32564 42484 32570
rect 42432 32506 42484 32512
rect 41696 32496 41748 32502
rect 41696 32438 41748 32444
rect 41512 32428 41564 32434
rect 41512 32370 41564 32376
rect 41880 32428 41932 32434
rect 41880 32370 41932 32376
rect 42248 32428 42300 32434
rect 42628 32416 42656 32710
rect 42708 32428 42760 32434
rect 42628 32388 42708 32416
rect 42248 32370 42300 32376
rect 42708 32370 42760 32376
rect 41420 32020 41472 32026
rect 41420 31962 41472 31968
rect 41512 31408 41564 31414
rect 41512 31350 41564 31356
rect 40960 31340 41012 31346
rect 40960 31282 41012 31288
rect 40592 30592 40644 30598
rect 40592 30534 40644 30540
rect 40500 30184 40552 30190
rect 40500 30126 40552 30132
rect 40500 30048 40552 30054
rect 40500 29990 40552 29996
rect 40408 29776 40460 29782
rect 40408 29718 40460 29724
rect 40420 29646 40448 29718
rect 40512 29714 40540 29990
rect 40500 29708 40552 29714
rect 40500 29650 40552 29656
rect 40408 29640 40460 29646
rect 40408 29582 40460 29588
rect 40604 29170 40632 30534
rect 40972 29646 41000 31282
rect 41328 30864 41380 30870
rect 41328 30806 41380 30812
rect 41340 30598 41368 30806
rect 41524 30802 41552 31350
rect 41512 30796 41564 30802
rect 41512 30738 41564 30744
rect 41328 30592 41380 30598
rect 41328 30534 41380 30540
rect 41524 30240 41552 30738
rect 41892 30326 41920 32370
rect 42260 31822 42288 32370
rect 42720 32026 42748 32370
rect 43076 32360 43128 32366
rect 43076 32302 43128 32308
rect 42708 32020 42760 32026
rect 42708 31962 42760 31968
rect 43088 31958 43116 32302
rect 43076 31952 43128 31958
rect 43076 31894 43128 31900
rect 42248 31816 42300 31822
rect 42248 31758 42300 31764
rect 41880 30320 41932 30326
rect 41880 30262 41932 30268
rect 41604 30252 41656 30258
rect 41524 30212 41604 30240
rect 40960 29640 41012 29646
rect 40960 29582 41012 29588
rect 41052 29504 41104 29510
rect 41052 29446 41104 29452
rect 40592 29164 40644 29170
rect 40592 29106 40644 29112
rect 40960 29164 41012 29170
rect 40960 29106 41012 29112
rect 40868 28960 40920 28966
rect 40868 28902 40920 28908
rect 40880 28762 40908 28902
rect 40868 28756 40920 28762
rect 40868 28698 40920 28704
rect 40776 28688 40828 28694
rect 40776 28630 40828 28636
rect 40788 28490 40816 28630
rect 40972 28558 41000 29106
rect 40960 28552 41012 28558
rect 40960 28494 41012 28500
rect 40684 28484 40736 28490
rect 40684 28426 40736 28432
rect 40776 28484 40828 28490
rect 40776 28426 40828 28432
rect 40696 28393 40724 28426
rect 40682 28384 40738 28393
rect 40682 28319 40738 28328
rect 40590 27432 40646 27441
rect 40590 27367 40646 27376
rect 40604 27334 40632 27367
rect 40592 27328 40644 27334
rect 40592 27270 40644 27276
rect 40500 27056 40552 27062
rect 40500 26998 40552 27004
rect 40408 26784 40460 26790
rect 40408 26726 40460 26732
rect 40316 26512 40368 26518
rect 40316 26454 40368 26460
rect 40316 25968 40368 25974
rect 40314 25936 40316 25945
rect 40368 25936 40370 25945
rect 40314 25871 40370 25880
rect 40316 25832 40368 25838
rect 40316 25774 40368 25780
rect 40328 25294 40356 25774
rect 40420 25702 40448 26726
rect 40512 26314 40540 26998
rect 40604 26382 40632 27270
rect 40696 26994 40724 28319
rect 40972 28150 41000 28494
rect 40960 28144 41012 28150
rect 40960 28086 41012 28092
rect 41064 27674 41092 29446
rect 41144 29028 41196 29034
rect 41144 28970 41196 28976
rect 41156 28558 41184 28970
rect 41144 28552 41196 28558
rect 41144 28494 41196 28500
rect 41052 27668 41104 27674
rect 41052 27610 41104 27616
rect 41064 26994 41092 27610
rect 40684 26988 40736 26994
rect 40684 26930 40736 26936
rect 41052 26988 41104 26994
rect 41052 26930 41104 26936
rect 40592 26376 40644 26382
rect 40592 26318 40644 26324
rect 40500 26308 40552 26314
rect 40500 26250 40552 26256
rect 40604 25906 40632 26318
rect 40868 26036 40920 26042
rect 40868 25978 40920 25984
rect 40880 25906 40908 25978
rect 40592 25900 40644 25906
rect 40592 25842 40644 25848
rect 40868 25900 40920 25906
rect 40868 25842 40920 25848
rect 40408 25696 40460 25702
rect 40408 25638 40460 25644
rect 40684 25696 40736 25702
rect 40684 25638 40736 25644
rect 40316 25288 40368 25294
rect 40316 25230 40368 25236
rect 40224 25152 40276 25158
rect 40224 25094 40276 25100
rect 40328 24970 40356 25230
rect 40236 24942 40356 24970
rect 40132 24608 40184 24614
rect 40132 24550 40184 24556
rect 40144 24206 40172 24550
rect 40236 24274 40264 24942
rect 40316 24744 40368 24750
rect 40316 24686 40368 24692
rect 40328 24410 40356 24686
rect 40316 24404 40368 24410
rect 40316 24346 40368 24352
rect 40224 24268 40276 24274
rect 40224 24210 40276 24216
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40040 23248 40092 23254
rect 40040 23190 40092 23196
rect 40420 23118 40448 25638
rect 40500 25288 40552 25294
rect 40500 25230 40552 25236
rect 40512 24886 40540 25230
rect 40500 24880 40552 24886
rect 40696 24857 40724 25638
rect 41156 25294 41184 28494
rect 41524 27470 41552 30212
rect 41604 30194 41656 30200
rect 42064 30184 42116 30190
rect 42064 30126 42116 30132
rect 42076 29646 42104 30126
rect 42260 29850 42288 31758
rect 43088 31482 43116 31894
rect 43076 31476 43128 31482
rect 43076 31418 43128 31424
rect 42432 30252 42484 30258
rect 42432 30194 42484 30200
rect 42708 30252 42760 30258
rect 42708 30194 42760 30200
rect 42248 29844 42300 29850
rect 42248 29786 42300 29792
rect 42064 29640 42116 29646
rect 42064 29582 42116 29588
rect 42444 29170 42472 30194
rect 42616 29708 42668 29714
rect 42616 29650 42668 29656
rect 42628 29306 42656 29650
rect 42720 29617 42748 30194
rect 42706 29608 42762 29617
rect 42706 29543 42762 29552
rect 43168 29572 43220 29578
rect 42616 29300 42668 29306
rect 42616 29242 42668 29248
rect 42720 29170 42748 29543
rect 43168 29514 43220 29520
rect 43180 29170 43208 29514
rect 42432 29164 42484 29170
rect 42432 29106 42484 29112
rect 42708 29164 42760 29170
rect 42708 29106 42760 29112
rect 43168 29164 43220 29170
rect 43168 29106 43220 29112
rect 42720 28994 42748 29106
rect 42720 28966 42932 28994
rect 42524 28960 42576 28966
rect 42524 28902 42576 28908
rect 42536 28694 42564 28902
rect 42524 28688 42576 28694
rect 42524 28630 42576 28636
rect 42904 28626 42932 28966
rect 42892 28620 42944 28626
rect 42892 28562 42944 28568
rect 41788 28552 41840 28558
rect 41788 28494 41840 28500
rect 41696 27668 41748 27674
rect 41696 27610 41748 27616
rect 41512 27464 41564 27470
rect 41512 27406 41564 27412
rect 41524 27130 41552 27406
rect 41708 27402 41736 27610
rect 41800 27470 41828 28494
rect 43272 28082 43300 34954
rect 43352 34604 43404 34610
rect 43456 34592 43484 35702
rect 43548 35698 43576 35974
rect 43536 35692 43588 35698
rect 43536 35634 43588 35640
rect 43628 35488 43680 35494
rect 43628 35430 43680 35436
rect 43640 35154 43668 35430
rect 43628 35148 43680 35154
rect 43628 35090 43680 35096
rect 43732 35018 43760 37828
rect 43904 35828 43956 35834
rect 43904 35770 43956 35776
rect 43720 35012 43772 35018
rect 43720 34954 43772 34960
rect 43916 34898 43944 35770
rect 43404 34564 43484 34592
rect 43824 34870 43944 34898
rect 43352 34546 43404 34552
rect 43364 34474 43392 34546
rect 43352 34468 43404 34474
rect 43352 34410 43404 34416
rect 43824 34134 43852 34870
rect 43904 34196 43956 34202
rect 43904 34138 43956 34144
rect 43812 34128 43864 34134
rect 43812 34070 43864 34076
rect 43916 33454 43944 34138
rect 43904 33448 43956 33454
rect 43904 33390 43956 33396
rect 43904 33312 43956 33318
rect 43902 33280 43904 33289
rect 43956 33280 43958 33289
rect 43902 33215 43958 33224
rect 43444 31816 43496 31822
rect 43444 31758 43496 31764
rect 43628 31816 43680 31822
rect 43628 31758 43680 31764
rect 43456 31210 43484 31758
rect 43640 31482 43668 31758
rect 44008 31754 44036 41386
rect 44192 39846 44220 43726
rect 44272 43104 44324 43110
rect 44272 43046 44324 43052
rect 44284 42838 44312 43046
rect 44272 42832 44324 42838
rect 44272 42774 44324 42780
rect 44376 42702 44404 44406
rect 44456 43240 44508 43246
rect 44456 43182 44508 43188
rect 44468 42770 44496 43182
rect 44456 42764 44508 42770
rect 44456 42706 44508 42712
rect 44364 42696 44416 42702
rect 44364 42638 44416 42644
rect 44180 39840 44232 39846
rect 44180 39782 44232 39788
rect 44364 39840 44416 39846
rect 44364 39782 44416 39788
rect 44088 39364 44140 39370
rect 44088 39306 44140 39312
rect 44100 38894 44128 39306
rect 44088 38888 44140 38894
rect 44088 38830 44140 38836
rect 44088 35692 44140 35698
rect 44088 35634 44140 35640
rect 44100 33114 44128 35634
rect 44192 35578 44220 39782
rect 44376 39642 44404 39782
rect 44364 39636 44416 39642
rect 44364 39578 44416 39584
rect 44364 38956 44416 38962
rect 44364 38898 44416 38904
rect 44272 38752 44324 38758
rect 44272 38694 44324 38700
rect 44284 36768 44312 38694
rect 44376 38486 44404 38898
rect 44456 38752 44508 38758
rect 44456 38694 44508 38700
rect 44364 38480 44416 38486
rect 44364 38422 44416 38428
rect 44468 38350 44496 38694
rect 44456 38344 44508 38350
rect 44456 38286 44508 38292
rect 44456 37120 44508 37126
rect 44456 37062 44508 37068
rect 44468 36786 44496 37062
rect 44456 36780 44508 36786
rect 44284 36740 44404 36768
rect 44272 36168 44324 36174
rect 44272 36110 44324 36116
rect 44284 35698 44312 36110
rect 44376 35834 44404 36740
rect 44456 36722 44508 36728
rect 44456 36032 44508 36038
rect 44456 35974 44508 35980
rect 44364 35828 44416 35834
rect 44364 35770 44416 35776
rect 44468 35698 44496 35974
rect 44272 35692 44324 35698
rect 44272 35634 44324 35640
rect 44456 35692 44508 35698
rect 44456 35634 44508 35640
rect 44364 35624 44416 35630
rect 44192 35550 44312 35578
rect 44364 35566 44416 35572
rect 44284 35193 44312 35550
rect 44270 35184 44326 35193
rect 44270 35119 44326 35128
rect 44284 35086 44312 35119
rect 44272 35080 44324 35086
rect 44272 35022 44324 35028
rect 44376 34746 44404 35566
rect 44468 34746 44496 35634
rect 44364 34740 44416 34746
rect 44364 34682 44416 34688
rect 44456 34740 44508 34746
rect 44456 34682 44508 34688
rect 44178 34640 44234 34649
rect 44456 34604 44508 34610
rect 44234 34584 44312 34592
rect 44178 34575 44180 34584
rect 44232 34564 44312 34584
rect 44180 34546 44232 34552
rect 44180 34400 44232 34406
rect 44180 34342 44232 34348
rect 44192 34066 44220 34342
rect 44284 34134 44312 34564
rect 44456 34546 44508 34552
rect 44272 34128 44324 34134
rect 44272 34070 44324 34076
rect 44180 34060 44232 34066
rect 44180 34002 44232 34008
rect 44364 33584 44416 33590
rect 44364 33526 44416 33532
rect 44180 33312 44232 33318
rect 44180 33254 44232 33260
rect 44192 33114 44220 33254
rect 44088 33108 44140 33114
rect 44088 33050 44140 33056
rect 44180 33108 44232 33114
rect 44180 33050 44232 33056
rect 44272 32768 44324 32774
rect 44272 32710 44324 32716
rect 44284 31822 44312 32710
rect 44272 31816 44324 31822
rect 44272 31758 44324 31764
rect 44008 31726 44128 31754
rect 43628 31476 43680 31482
rect 43628 31418 43680 31424
rect 43536 31340 43588 31346
rect 43536 31282 43588 31288
rect 43444 31204 43496 31210
rect 43444 31146 43496 31152
rect 43548 31090 43576 31282
rect 43456 31062 43576 31090
rect 43456 30734 43484 31062
rect 43444 30728 43496 30734
rect 43444 30670 43496 30676
rect 43456 30394 43484 30670
rect 43536 30592 43588 30598
rect 43536 30534 43588 30540
rect 43444 30388 43496 30394
rect 43444 30330 43496 30336
rect 43548 30326 43576 30534
rect 43536 30320 43588 30326
rect 43536 30262 43588 30268
rect 43996 30252 44048 30258
rect 43996 30194 44048 30200
rect 43352 30184 43404 30190
rect 43352 30126 43404 30132
rect 43812 30184 43864 30190
rect 43812 30126 43864 30132
rect 43364 29306 43392 30126
rect 43536 30116 43588 30122
rect 43536 30058 43588 30064
rect 43548 29782 43576 30058
rect 43536 29776 43588 29782
rect 43536 29718 43588 29724
rect 43444 29708 43496 29714
rect 43444 29650 43496 29656
rect 43352 29300 43404 29306
rect 43352 29242 43404 29248
rect 43456 29238 43484 29650
rect 43548 29510 43576 29718
rect 43824 29646 43852 30126
rect 44008 29646 44036 30194
rect 43812 29640 43864 29646
rect 43718 29608 43774 29617
rect 43812 29582 43864 29588
rect 43996 29640 44048 29646
rect 43996 29582 44048 29588
rect 43718 29543 43720 29552
rect 43772 29543 43774 29552
rect 43720 29514 43772 29520
rect 43536 29504 43588 29510
rect 43536 29446 43588 29452
rect 43444 29232 43496 29238
rect 43444 29174 43496 29180
rect 43352 28620 43404 28626
rect 43352 28562 43404 28568
rect 43364 28218 43392 28562
rect 43352 28212 43404 28218
rect 43352 28154 43404 28160
rect 43444 28144 43496 28150
rect 43444 28086 43496 28092
rect 43260 28076 43312 28082
rect 43260 28018 43312 28024
rect 41788 27464 41840 27470
rect 42340 27464 42392 27470
rect 41788 27406 41840 27412
rect 42338 27432 42340 27441
rect 42392 27432 42394 27441
rect 41696 27396 41748 27402
rect 41696 27338 41748 27344
rect 41512 27124 41564 27130
rect 41512 27066 41564 27072
rect 41236 27056 41288 27062
rect 41236 26998 41288 27004
rect 41248 25294 41276 26998
rect 41800 26382 41828 27406
rect 43272 27402 43300 28018
rect 42338 27367 42394 27376
rect 42800 27396 42852 27402
rect 42800 27338 42852 27344
rect 43260 27396 43312 27402
rect 43260 27338 43312 27344
rect 42340 27328 42392 27334
rect 42340 27270 42392 27276
rect 42352 27062 42380 27270
rect 42340 27056 42392 27062
rect 42340 26998 42392 27004
rect 42812 26994 42840 27338
rect 42800 26988 42852 26994
rect 42800 26930 42852 26936
rect 43456 26518 43484 28086
rect 43548 26926 43576 29446
rect 44008 29102 44036 29582
rect 43996 29096 44048 29102
rect 43996 29038 44048 29044
rect 43720 28552 43772 28558
rect 43720 28494 43772 28500
rect 43732 27674 43760 28494
rect 43904 28416 43956 28422
rect 43904 28358 43956 28364
rect 43916 28014 43944 28358
rect 43904 28008 43956 28014
rect 43904 27950 43956 27956
rect 43812 27872 43864 27878
rect 43812 27814 43864 27820
rect 43904 27872 43956 27878
rect 43904 27814 43956 27820
rect 43720 27668 43772 27674
rect 43720 27610 43772 27616
rect 43720 26988 43772 26994
rect 43720 26930 43772 26936
rect 43536 26920 43588 26926
rect 43536 26862 43588 26868
rect 43444 26512 43496 26518
rect 43496 26472 43576 26500
rect 43444 26454 43496 26460
rect 41420 26376 41472 26382
rect 41420 26318 41472 26324
rect 41604 26376 41656 26382
rect 41604 26318 41656 26324
rect 41788 26376 41840 26382
rect 41788 26318 41840 26324
rect 43076 26376 43128 26382
rect 43076 26318 43128 26324
rect 41432 25838 41460 26318
rect 41616 25906 41644 26318
rect 41880 26308 41932 26314
rect 41880 26250 41932 26256
rect 41696 26240 41748 26246
rect 41696 26182 41748 26188
rect 41604 25900 41656 25906
rect 41604 25842 41656 25848
rect 41420 25832 41472 25838
rect 41420 25774 41472 25780
rect 41708 25702 41736 26182
rect 41788 25900 41840 25906
rect 41788 25842 41840 25848
rect 41696 25696 41748 25702
rect 41696 25638 41748 25644
rect 41144 25288 41196 25294
rect 41144 25230 41196 25236
rect 41236 25288 41288 25294
rect 41236 25230 41288 25236
rect 40960 25220 41012 25226
rect 40960 25162 41012 25168
rect 40500 24822 40552 24828
rect 40682 24848 40738 24857
rect 40682 24783 40738 24792
rect 40408 23112 40460 23118
rect 40408 23054 40460 23060
rect 40696 22982 40724 24783
rect 40972 24682 41000 25162
rect 41248 24886 41276 25230
rect 41420 25152 41472 25158
rect 41420 25094 41472 25100
rect 41432 24954 41460 25094
rect 41420 24948 41472 24954
rect 41420 24890 41472 24896
rect 41236 24880 41288 24886
rect 41236 24822 41288 24828
rect 41052 24812 41104 24818
rect 41052 24754 41104 24760
rect 40960 24676 41012 24682
rect 40960 24618 41012 24624
rect 41064 24070 41092 24754
rect 41248 24138 41276 24822
rect 41432 24818 41460 24890
rect 41420 24812 41472 24818
rect 41420 24754 41472 24760
rect 41708 24206 41736 25638
rect 41800 25158 41828 25842
rect 41788 25152 41840 25158
rect 41788 25094 41840 25100
rect 41892 24750 41920 26250
rect 42800 26240 42852 26246
rect 42800 26182 42852 26188
rect 42812 25650 42840 26182
rect 42720 25622 43024 25650
rect 42720 25294 42748 25622
rect 42800 25492 42852 25498
rect 42800 25434 42852 25440
rect 42708 25288 42760 25294
rect 42708 25230 42760 25236
rect 41972 25220 42024 25226
rect 41972 25162 42024 25168
rect 41880 24744 41932 24750
rect 41880 24686 41932 24692
rect 41892 24206 41920 24686
rect 41984 24342 42012 25162
rect 42812 24682 42840 25434
rect 42892 25288 42944 25294
rect 42892 25230 42944 25236
rect 42904 24954 42932 25230
rect 42892 24948 42944 24954
rect 42892 24890 42944 24896
rect 42996 24818 43024 25622
rect 43088 25294 43116 26318
rect 43548 25906 43576 26472
rect 43732 26450 43760 26930
rect 43720 26444 43772 26450
rect 43720 26386 43772 26392
rect 43732 26042 43760 26386
rect 43824 26314 43852 27814
rect 43916 27470 43944 27814
rect 43904 27464 43956 27470
rect 43904 27406 43956 27412
rect 43812 26308 43864 26314
rect 43812 26250 43864 26256
rect 43720 26036 43772 26042
rect 43720 25978 43772 25984
rect 43444 25900 43496 25906
rect 43444 25842 43496 25848
rect 43536 25900 43588 25906
rect 43536 25842 43588 25848
rect 43456 25294 43484 25842
rect 43076 25288 43128 25294
rect 43076 25230 43128 25236
rect 43444 25288 43496 25294
rect 43444 25230 43496 25236
rect 42984 24812 43036 24818
rect 42984 24754 43036 24760
rect 42800 24676 42852 24682
rect 42800 24618 42852 24624
rect 41972 24336 42024 24342
rect 41972 24278 42024 24284
rect 42800 24336 42852 24342
rect 42800 24278 42852 24284
rect 42812 24206 42840 24278
rect 42996 24206 43024 24754
rect 43456 24614 43484 25230
rect 43626 24712 43682 24721
rect 43626 24647 43628 24656
rect 43680 24647 43682 24656
rect 43628 24618 43680 24624
rect 43444 24608 43496 24614
rect 43444 24550 43496 24556
rect 43076 24336 43128 24342
rect 43076 24278 43128 24284
rect 41696 24200 41748 24206
rect 41696 24142 41748 24148
rect 41880 24200 41932 24206
rect 41880 24142 41932 24148
rect 42800 24200 42852 24206
rect 42800 24142 42852 24148
rect 42984 24200 43036 24206
rect 42984 24142 43036 24148
rect 41236 24132 41288 24138
rect 41236 24074 41288 24080
rect 42892 24132 42944 24138
rect 42892 24074 42944 24080
rect 41052 24064 41104 24070
rect 41052 24006 41104 24012
rect 42904 23118 42932 24074
rect 43088 23118 43116 24278
rect 43640 24138 43668 24618
rect 43628 24132 43680 24138
rect 43628 24074 43680 24080
rect 43260 23792 43312 23798
rect 43260 23734 43312 23740
rect 43272 23186 43300 23734
rect 43824 23730 43852 26250
rect 43352 23724 43404 23730
rect 43352 23666 43404 23672
rect 43812 23724 43864 23730
rect 43812 23666 43864 23672
rect 43260 23180 43312 23186
rect 43260 23122 43312 23128
rect 42892 23112 42944 23118
rect 42892 23054 42944 23060
rect 43076 23112 43128 23118
rect 43076 23054 43128 23060
rect 40684 22976 40736 22982
rect 40684 22918 40736 22924
rect 43272 22642 43300 23122
rect 43364 22982 43392 23666
rect 43720 23044 43772 23050
rect 43720 22986 43772 22992
rect 43352 22976 43404 22982
rect 43352 22918 43404 22924
rect 43536 22976 43588 22982
rect 43536 22918 43588 22924
rect 43548 22642 43576 22918
rect 43732 22778 43760 22986
rect 43720 22772 43772 22778
rect 43720 22714 43772 22720
rect 43260 22636 43312 22642
rect 43260 22578 43312 22584
rect 43536 22636 43588 22642
rect 43536 22578 43588 22584
rect 43272 22234 43300 22578
rect 43260 22228 43312 22234
rect 43260 22170 43312 22176
rect 43548 21962 43576 22578
rect 43824 22098 43852 23666
rect 43916 23322 43944 27406
rect 44100 26874 44128 31726
rect 44284 31278 44312 31758
rect 44272 31272 44324 31278
rect 44272 31214 44324 31220
rect 44376 31142 44404 33526
rect 44468 32978 44496 34546
rect 44456 32972 44508 32978
rect 44456 32914 44508 32920
rect 44456 32428 44508 32434
rect 44456 32370 44508 32376
rect 44468 32298 44496 32370
rect 44456 32292 44508 32298
rect 44456 32234 44508 32240
rect 44468 31822 44496 32234
rect 44456 31816 44508 31822
rect 44456 31758 44508 31764
rect 44560 31754 44588 45834
rect 44824 44396 44876 44402
rect 44824 44338 44876 44344
rect 44836 43994 44864 44338
rect 44824 43988 44876 43994
rect 44824 43930 44876 43936
rect 44928 43858 44956 45902
rect 45664 45830 45692 47602
rect 45848 47569 45876 48010
rect 46204 48000 46256 48006
rect 46204 47942 46256 47948
rect 46112 47796 46164 47802
rect 46112 47738 46164 47744
rect 46124 47598 46152 47738
rect 46216 47666 46244 47942
rect 46204 47660 46256 47666
rect 46204 47602 46256 47608
rect 46112 47592 46164 47598
rect 45834 47560 45890 47569
rect 46112 47534 46164 47540
rect 45834 47495 45890 47504
rect 45744 46980 45796 46986
rect 45744 46922 45796 46928
rect 45756 46578 45784 46922
rect 45744 46572 45796 46578
rect 45744 46514 45796 46520
rect 45756 46170 45784 46514
rect 45744 46164 45796 46170
rect 45744 46106 45796 46112
rect 45008 45824 45060 45830
rect 45008 45766 45060 45772
rect 45652 45824 45704 45830
rect 45652 45766 45704 45772
rect 44916 43852 44968 43858
rect 44916 43794 44968 43800
rect 44916 43716 44968 43722
rect 44916 43658 44968 43664
rect 44638 43480 44694 43489
rect 44638 43415 44640 43424
rect 44692 43415 44694 43424
rect 44640 43386 44692 43392
rect 44928 43382 44956 43658
rect 44916 43376 44968 43382
rect 44916 43318 44968 43324
rect 45020 43314 45048 45766
rect 45848 45558 45876 47495
rect 45928 47456 45980 47462
rect 45928 47398 45980 47404
rect 46112 47456 46164 47462
rect 46112 47398 46164 47404
rect 45940 47054 45968 47398
rect 45928 47048 45980 47054
rect 45928 46990 45980 46996
rect 45836 45552 45888 45558
rect 45836 45494 45888 45500
rect 45928 45484 45980 45490
rect 45928 45426 45980 45432
rect 45376 45280 45428 45286
rect 45376 45222 45428 45228
rect 45744 45280 45796 45286
rect 45744 45222 45796 45228
rect 45190 44160 45246 44169
rect 45190 44095 45246 44104
rect 45204 43858 45232 44095
rect 45192 43852 45244 43858
rect 45244 43812 45324 43840
rect 45192 43794 45244 43800
rect 45008 43308 45060 43314
rect 45008 43250 45060 43256
rect 45020 42702 45048 43250
rect 45192 43240 45244 43246
rect 45192 43182 45244 43188
rect 45204 42702 45232 43182
rect 45008 42696 45060 42702
rect 45006 42664 45008 42673
rect 45192 42696 45244 42702
rect 45060 42664 45062 42673
rect 45192 42638 45244 42644
rect 45006 42599 45062 42608
rect 45192 42560 45244 42566
rect 45192 42502 45244 42508
rect 45204 41614 45232 42502
rect 45192 41608 45244 41614
rect 45192 41550 45244 41556
rect 45204 40458 45232 41550
rect 45296 41478 45324 43812
rect 45388 43722 45416 45222
rect 45560 44736 45612 44742
rect 45560 44678 45612 44684
rect 45468 44396 45520 44402
rect 45468 44338 45520 44344
rect 45376 43716 45428 43722
rect 45376 43658 45428 43664
rect 45480 43314 45508 44338
rect 45572 43926 45600 44678
rect 45560 43920 45612 43926
rect 45560 43862 45612 43868
rect 45650 43888 45706 43897
rect 45572 43704 45600 43862
rect 45756 43858 45784 45222
rect 45834 44296 45890 44305
rect 45834 44231 45836 44240
rect 45888 44231 45890 44240
rect 45836 44202 45888 44208
rect 45650 43823 45652 43832
rect 45704 43823 45706 43832
rect 45744 43852 45796 43858
rect 45652 43794 45704 43800
rect 45744 43794 45796 43800
rect 45652 43716 45704 43722
rect 45572 43676 45652 43704
rect 45652 43658 45704 43664
rect 45560 43444 45612 43450
rect 45560 43386 45612 43392
rect 45572 43314 45600 43386
rect 45468 43308 45520 43314
rect 45468 43250 45520 43256
rect 45560 43308 45612 43314
rect 45560 43250 45612 43256
rect 45836 43308 45888 43314
rect 45836 43250 45888 43256
rect 45376 42900 45428 42906
rect 45376 42842 45428 42848
rect 45388 42702 45416 42842
rect 45376 42696 45428 42702
rect 45376 42638 45428 42644
rect 45560 42696 45612 42702
rect 45560 42638 45612 42644
rect 45572 41682 45600 42638
rect 45560 41676 45612 41682
rect 45560 41618 45612 41624
rect 45284 41472 45336 41478
rect 45336 41432 45508 41460
rect 45284 41414 45336 41420
rect 45192 40452 45244 40458
rect 45192 40394 45244 40400
rect 44824 40044 44876 40050
rect 44824 39986 44876 39992
rect 44836 39370 44864 39986
rect 45100 39840 45152 39846
rect 45100 39782 45152 39788
rect 45008 39568 45060 39574
rect 45008 39510 45060 39516
rect 45020 39438 45048 39510
rect 45008 39432 45060 39438
rect 45008 39374 45060 39380
rect 44824 39364 44876 39370
rect 44824 39306 44876 39312
rect 44732 39296 44784 39302
rect 44732 39238 44784 39244
rect 44744 38962 44772 39238
rect 45020 38962 45048 39374
rect 45112 39302 45140 39782
rect 45204 39642 45232 40394
rect 45376 39840 45428 39846
rect 45376 39782 45428 39788
rect 45192 39636 45244 39642
rect 45192 39578 45244 39584
rect 45284 39636 45336 39642
rect 45284 39578 45336 39584
rect 45296 39438 45324 39578
rect 45284 39432 45336 39438
rect 45284 39374 45336 39380
rect 45192 39364 45244 39370
rect 45192 39306 45244 39312
rect 45100 39296 45152 39302
rect 45100 39238 45152 39244
rect 44732 38956 44784 38962
rect 44732 38898 44784 38904
rect 45008 38956 45060 38962
rect 45008 38898 45060 38904
rect 44732 38820 44784 38826
rect 44732 38762 44784 38768
rect 44640 38752 44692 38758
rect 44640 38694 44692 38700
rect 44652 36582 44680 38694
rect 44744 38554 44772 38762
rect 44732 38548 44784 38554
rect 44732 38490 44784 38496
rect 45204 38418 45232 39306
rect 45192 38412 45244 38418
rect 45192 38354 45244 38360
rect 44824 38208 44876 38214
rect 44824 38150 44876 38156
rect 44732 37800 44784 37806
rect 44732 37742 44784 37748
rect 44744 37466 44772 37742
rect 44732 37460 44784 37466
rect 44732 37402 44784 37408
rect 44744 37330 44772 37402
rect 44732 37324 44784 37330
rect 44732 37266 44784 37272
rect 44836 36922 44864 38150
rect 45204 37466 45232 38354
rect 45296 38049 45324 39374
rect 45388 39030 45416 39782
rect 45376 39024 45428 39030
rect 45376 38966 45428 38972
rect 45480 38962 45508 41432
rect 45848 40118 45876 43250
rect 45940 43110 45968 45426
rect 46124 44198 46152 47398
rect 46216 46510 46244 47602
rect 46308 47530 46336 48078
rect 46388 48068 46440 48074
rect 46388 48010 46440 48016
rect 46296 47524 46348 47530
rect 46296 47466 46348 47472
rect 46400 46918 46428 48010
rect 46584 47666 46612 48146
rect 47400 48136 47452 48142
rect 47400 48078 47452 48084
rect 46940 48068 46992 48074
rect 46940 48010 46992 48016
rect 46952 47802 46980 48010
rect 46940 47796 46992 47802
rect 46940 47738 46992 47744
rect 46572 47660 46624 47666
rect 46572 47602 46624 47608
rect 46584 47462 46612 47602
rect 46572 47456 46624 47462
rect 46572 47398 46624 47404
rect 46952 47054 46980 47738
rect 47032 47592 47084 47598
rect 47032 47534 47084 47540
rect 46940 47048 46992 47054
rect 46940 46990 46992 46996
rect 46388 46912 46440 46918
rect 46388 46854 46440 46860
rect 46848 46572 46900 46578
rect 46848 46514 46900 46520
rect 46204 46504 46256 46510
rect 46204 46446 46256 46452
rect 46296 45892 46348 45898
rect 46296 45834 46348 45840
rect 46112 44192 46164 44198
rect 46112 44134 46164 44140
rect 46020 43988 46072 43994
rect 46020 43930 46072 43936
rect 46032 43625 46060 43930
rect 46204 43648 46256 43654
rect 46018 43616 46074 43625
rect 46204 43590 46256 43596
rect 46018 43551 46074 43560
rect 46216 43450 46244 43590
rect 46204 43444 46256 43450
rect 46204 43386 46256 43392
rect 45928 43104 45980 43110
rect 45928 43046 45980 43052
rect 46308 41138 46336 45834
rect 46480 45484 46532 45490
rect 46480 45426 46532 45432
rect 46492 44878 46520 45426
rect 46860 45422 46888 46514
rect 46848 45416 46900 45422
rect 46848 45358 46900 45364
rect 46572 45076 46624 45082
rect 46572 45018 46624 45024
rect 46480 44872 46532 44878
rect 46480 44814 46532 44820
rect 46492 43874 46520 44814
rect 46584 44334 46612 45018
rect 47044 44878 47072 47534
rect 47124 47048 47176 47054
rect 47124 46990 47176 46996
rect 47216 47048 47268 47054
rect 47216 46990 47268 46996
rect 47136 45898 47164 46990
rect 47124 45892 47176 45898
rect 47124 45834 47176 45840
rect 47136 45490 47164 45834
rect 47228 45830 47256 46990
rect 47216 45824 47268 45830
rect 47216 45766 47268 45772
rect 47124 45484 47176 45490
rect 47124 45426 47176 45432
rect 47136 45082 47164 45426
rect 47216 45348 47268 45354
rect 47216 45290 47268 45296
rect 47124 45076 47176 45082
rect 47124 45018 47176 45024
rect 47032 44872 47084 44878
rect 47032 44814 47084 44820
rect 46664 44396 46716 44402
rect 46664 44338 46716 44344
rect 46572 44328 46624 44334
rect 46676 44305 46704 44338
rect 46572 44270 46624 44276
rect 46662 44296 46718 44305
rect 46584 44169 46612 44270
rect 46662 44231 46718 44240
rect 46570 44160 46626 44169
rect 46570 44095 46626 44104
rect 46848 43920 46900 43926
rect 46492 43846 46612 43874
rect 46848 43862 46900 43868
rect 46480 43784 46532 43790
rect 46480 43726 46532 43732
rect 46492 43450 46520 43726
rect 46480 43444 46532 43450
rect 46480 43386 46532 43392
rect 46584 43314 46612 43846
rect 46756 43852 46808 43858
rect 46756 43794 46808 43800
rect 46572 43308 46624 43314
rect 46572 43250 46624 43256
rect 46388 43240 46440 43246
rect 46388 43182 46440 43188
rect 46400 42906 46428 43182
rect 46480 43104 46532 43110
rect 46480 43046 46532 43052
rect 46388 42900 46440 42906
rect 46388 42842 46440 42848
rect 46492 42634 46520 43046
rect 46584 42702 46612 43250
rect 46768 42906 46796 43794
rect 46756 42900 46808 42906
rect 46756 42842 46808 42848
rect 46572 42696 46624 42702
rect 46572 42638 46624 42644
rect 46480 42628 46532 42634
rect 46480 42570 46532 42576
rect 46492 42158 46520 42570
rect 46480 42152 46532 42158
rect 46480 42094 46532 42100
rect 45928 41132 45980 41138
rect 45928 41074 45980 41080
rect 46296 41132 46348 41138
rect 46296 41074 46348 41080
rect 45560 40112 45612 40118
rect 45560 40054 45612 40060
rect 45836 40112 45888 40118
rect 45836 40054 45888 40060
rect 45572 39982 45600 40054
rect 45560 39976 45612 39982
rect 45560 39918 45612 39924
rect 45560 39840 45612 39846
rect 45560 39782 45612 39788
rect 45572 39574 45600 39782
rect 45560 39568 45612 39574
rect 45560 39510 45612 39516
rect 45652 39432 45704 39438
rect 45652 39374 45704 39380
rect 45664 39098 45692 39374
rect 45652 39092 45704 39098
rect 45652 39034 45704 39040
rect 45468 38956 45520 38962
rect 45468 38898 45520 38904
rect 45836 38956 45888 38962
rect 45836 38898 45888 38904
rect 45560 38888 45612 38894
rect 45560 38830 45612 38836
rect 45282 38040 45338 38049
rect 45282 37975 45338 37984
rect 45376 38004 45428 38010
rect 45376 37946 45428 37952
rect 45192 37460 45244 37466
rect 45192 37402 45244 37408
rect 45388 37330 45416 37946
rect 45572 37874 45600 38830
rect 45744 38752 45796 38758
rect 45664 38712 45744 38740
rect 45560 37868 45612 37874
rect 45560 37810 45612 37816
rect 45376 37324 45428 37330
rect 45376 37266 45428 37272
rect 45284 37256 45336 37262
rect 45284 37198 45336 37204
rect 44824 36916 44876 36922
rect 44824 36858 44876 36864
rect 44640 36576 44692 36582
rect 44640 36518 44692 36524
rect 45296 36174 45324 37198
rect 45572 36378 45600 37810
rect 45664 37738 45692 38712
rect 45744 38694 45796 38700
rect 45848 37806 45876 38898
rect 45836 37800 45888 37806
rect 45836 37742 45888 37748
rect 45652 37732 45704 37738
rect 45652 37674 45704 37680
rect 45652 37120 45704 37126
rect 45652 37062 45704 37068
rect 45560 36372 45612 36378
rect 45560 36314 45612 36320
rect 45284 36168 45336 36174
rect 45284 36110 45336 36116
rect 45192 35760 45244 35766
rect 45192 35702 45244 35708
rect 45008 35692 45060 35698
rect 45008 35634 45060 35640
rect 45020 35086 45048 35634
rect 45100 35488 45152 35494
rect 45100 35430 45152 35436
rect 45112 35154 45140 35430
rect 45100 35148 45152 35154
rect 45100 35090 45152 35096
rect 45008 35080 45060 35086
rect 45008 35022 45060 35028
rect 44916 35012 44968 35018
rect 44916 34954 44968 34960
rect 44824 34536 44876 34542
rect 44824 34478 44876 34484
rect 44732 34400 44784 34406
rect 44732 34342 44784 34348
rect 44640 33312 44692 33318
rect 44744 33300 44772 34342
rect 44692 33272 44772 33300
rect 44640 33254 44692 33260
rect 44836 32910 44864 34478
rect 44928 34082 44956 34954
rect 45204 34610 45232 35702
rect 45100 34604 45152 34610
rect 45100 34546 45152 34552
rect 45192 34604 45244 34610
rect 45192 34546 45244 34552
rect 45008 34400 45060 34406
rect 45008 34342 45060 34348
rect 45020 34202 45048 34342
rect 45008 34196 45060 34202
rect 45008 34138 45060 34144
rect 44928 34054 45048 34082
rect 44916 33992 44968 33998
rect 44916 33934 44968 33940
rect 44928 33674 44956 33934
rect 45020 33930 45048 34054
rect 45112 33998 45140 34546
rect 45204 34474 45232 34546
rect 45192 34468 45244 34474
rect 45192 34410 45244 34416
rect 45100 33992 45152 33998
rect 45100 33934 45152 33940
rect 45008 33924 45060 33930
rect 45008 33866 45060 33872
rect 44928 33646 45140 33674
rect 45204 33658 45232 34410
rect 45112 33590 45140 33646
rect 45192 33652 45244 33658
rect 45192 33594 45244 33600
rect 45100 33584 45152 33590
rect 45100 33526 45152 33532
rect 44916 33516 44968 33522
rect 44916 33458 44968 33464
rect 44928 33114 44956 33458
rect 44916 33108 44968 33114
rect 44916 33050 44968 33056
rect 44824 32904 44876 32910
rect 44824 32846 44876 32852
rect 44824 32224 44876 32230
rect 44824 32166 44876 32172
rect 44560 31726 44680 31754
rect 44456 31272 44508 31278
rect 44456 31214 44508 31220
rect 44180 31136 44232 31142
rect 44180 31078 44232 31084
rect 44364 31136 44416 31142
rect 44364 31078 44416 31084
rect 44192 29646 44220 31078
rect 44272 30728 44324 30734
rect 44272 30670 44324 30676
rect 44180 29640 44232 29646
rect 44180 29582 44232 29588
rect 44192 29170 44220 29582
rect 44284 29306 44312 30670
rect 44364 30660 44416 30666
rect 44364 30602 44416 30608
rect 44272 29300 44324 29306
rect 44272 29242 44324 29248
rect 44180 29164 44232 29170
rect 44180 29106 44232 29112
rect 44376 28218 44404 30602
rect 44364 28212 44416 28218
rect 44364 28154 44416 28160
rect 44008 26846 44128 26874
rect 44008 26246 44036 26846
rect 44088 26784 44140 26790
rect 44088 26726 44140 26732
rect 43996 26240 44048 26246
rect 43996 26182 44048 26188
rect 44100 25770 44128 26726
rect 44468 26518 44496 31214
rect 44548 30796 44600 30802
rect 44548 30738 44600 30744
rect 44560 30394 44588 30738
rect 44548 30388 44600 30394
rect 44548 30330 44600 30336
rect 44652 27130 44680 31726
rect 44836 31346 44864 32166
rect 44824 31340 44876 31346
rect 44824 31282 44876 31288
rect 44732 31136 44784 31142
rect 44732 31078 44784 31084
rect 44744 30666 44772 31078
rect 44836 30938 44864 31282
rect 44824 30932 44876 30938
rect 44824 30874 44876 30880
rect 44732 30660 44784 30666
rect 44732 30602 44784 30608
rect 44928 30326 44956 33050
rect 45296 32910 45324 36110
rect 45468 36100 45520 36106
rect 45468 36042 45520 36048
rect 45480 35222 45508 36042
rect 45468 35216 45520 35222
rect 45664 35204 45692 37062
rect 45848 36786 45876 37742
rect 45836 36780 45888 36786
rect 45836 36722 45888 36728
rect 45468 35158 45520 35164
rect 45572 35176 45692 35204
rect 45480 34542 45508 35158
rect 45468 34536 45520 34542
rect 45468 34478 45520 34484
rect 45376 33924 45428 33930
rect 45376 33866 45428 33872
rect 45388 33114 45416 33866
rect 45572 33658 45600 35176
rect 45940 35018 45968 41074
rect 46860 40594 46888 43862
rect 46940 43444 46992 43450
rect 46940 43386 46992 43392
rect 46952 43110 46980 43386
rect 46940 43104 46992 43110
rect 46940 43046 46992 43052
rect 46940 40928 46992 40934
rect 46940 40870 46992 40876
rect 46848 40588 46900 40594
rect 46848 40530 46900 40536
rect 46664 40520 46716 40526
rect 46664 40462 46716 40468
rect 46480 40452 46532 40458
rect 46480 40394 46532 40400
rect 46572 40452 46624 40458
rect 46572 40394 46624 40400
rect 46492 39846 46520 40394
rect 46584 40050 46612 40394
rect 46676 40118 46704 40462
rect 46952 40186 46980 40870
rect 46940 40180 46992 40186
rect 46940 40122 46992 40128
rect 46664 40112 46716 40118
rect 46664 40054 46716 40060
rect 46572 40044 46624 40050
rect 46572 39986 46624 39992
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46676 39574 46704 40054
rect 46664 39568 46716 39574
rect 46664 39510 46716 39516
rect 46020 39092 46072 39098
rect 46020 39034 46072 39040
rect 46032 38350 46060 39034
rect 46952 38894 46980 40122
rect 46940 38888 46992 38894
rect 46940 38830 46992 38836
rect 46296 38820 46348 38826
rect 46296 38762 46348 38768
rect 46308 38554 46336 38762
rect 46940 38752 46992 38758
rect 46940 38694 46992 38700
rect 46386 38584 46442 38593
rect 46112 38548 46164 38554
rect 46112 38490 46164 38496
rect 46296 38548 46348 38554
rect 46386 38519 46442 38528
rect 46296 38490 46348 38496
rect 46020 38344 46072 38350
rect 46020 38286 46072 38292
rect 46032 37466 46060 38286
rect 46124 37874 46152 38490
rect 46400 38486 46428 38519
rect 46204 38480 46256 38486
rect 46204 38422 46256 38428
rect 46388 38480 46440 38486
rect 46388 38422 46440 38428
rect 46216 38214 46244 38422
rect 46952 38350 46980 38694
rect 46388 38344 46440 38350
rect 46756 38344 46808 38350
rect 46440 38328 46704 38332
rect 46440 38322 46716 38328
rect 46440 38304 46664 38322
rect 46388 38286 46440 38292
rect 46296 38276 46348 38282
rect 46756 38286 46808 38292
rect 46940 38344 46992 38350
rect 46940 38286 46992 38292
rect 46664 38264 46716 38270
rect 46296 38218 46348 38224
rect 46204 38208 46256 38214
rect 46204 38150 46256 38156
rect 46112 37868 46164 37874
rect 46112 37810 46164 37816
rect 46020 37460 46072 37466
rect 46020 37402 46072 37408
rect 46124 37262 46152 37810
rect 46216 37806 46244 38150
rect 46204 37800 46256 37806
rect 46204 37742 46256 37748
rect 46308 37330 46336 38218
rect 46768 38010 46796 38286
rect 46756 38004 46808 38010
rect 46756 37946 46808 37952
rect 46480 37868 46532 37874
rect 46480 37810 46532 37816
rect 46388 37800 46440 37806
rect 46388 37742 46440 37748
rect 46400 37398 46428 37742
rect 46388 37392 46440 37398
rect 46388 37334 46440 37340
rect 46296 37324 46348 37330
rect 46296 37266 46348 37272
rect 46492 37262 46520 37810
rect 46112 37256 46164 37262
rect 46112 37198 46164 37204
rect 46204 37256 46256 37262
rect 46204 37198 46256 37204
rect 46480 37256 46532 37262
rect 46480 37198 46532 37204
rect 46124 36174 46152 37198
rect 46216 36174 46244 37198
rect 46756 36780 46808 36786
rect 46756 36722 46808 36728
rect 46112 36168 46164 36174
rect 46112 36110 46164 36116
rect 46204 36168 46256 36174
rect 46204 36110 46256 36116
rect 46124 35630 46152 36110
rect 46216 35834 46244 36110
rect 46204 35828 46256 35834
rect 46204 35770 46256 35776
rect 46296 35760 46348 35766
rect 46296 35702 46348 35708
rect 46112 35624 46164 35630
rect 46112 35566 46164 35572
rect 45928 35012 45980 35018
rect 45928 34954 45980 34960
rect 46308 34950 46336 35702
rect 46388 35692 46440 35698
rect 46388 35634 46440 35640
rect 46400 35086 46428 35634
rect 46388 35080 46440 35086
rect 46388 35022 46440 35028
rect 46296 34944 46348 34950
rect 46296 34886 46348 34892
rect 45742 34504 45798 34513
rect 45742 34439 45798 34448
rect 45756 34134 45784 34439
rect 46308 34202 46336 34886
rect 46296 34196 46348 34202
rect 46296 34138 46348 34144
rect 45744 34128 45796 34134
rect 45744 34070 45796 34076
rect 45560 33652 45612 33658
rect 45560 33594 45612 33600
rect 45560 33312 45612 33318
rect 45480 33260 45560 33266
rect 45480 33254 45612 33260
rect 45480 33238 45600 33254
rect 45376 33108 45428 33114
rect 45376 33050 45428 33056
rect 45284 32904 45336 32910
rect 45284 32846 45336 32852
rect 45192 32768 45244 32774
rect 45192 32710 45244 32716
rect 45204 32434 45232 32710
rect 45008 32428 45060 32434
rect 45008 32370 45060 32376
rect 45192 32428 45244 32434
rect 45192 32370 45244 32376
rect 45020 31822 45048 32370
rect 45204 31890 45232 32370
rect 45192 31884 45244 31890
rect 45192 31826 45244 31832
rect 45008 31816 45060 31822
rect 45008 31758 45060 31764
rect 45284 31476 45336 31482
rect 45284 31418 45336 31424
rect 45296 31278 45324 31418
rect 45284 31272 45336 31278
rect 45284 31214 45336 31220
rect 45296 30802 45324 31214
rect 45284 30796 45336 30802
rect 45284 30738 45336 30744
rect 45480 30394 45508 33238
rect 46112 31340 46164 31346
rect 46112 31282 46164 31288
rect 45468 30388 45520 30394
rect 45468 30330 45520 30336
rect 44916 30320 44968 30326
rect 44916 30262 44968 30268
rect 45192 30252 45244 30258
rect 45192 30194 45244 30200
rect 44916 30184 44968 30190
rect 44916 30126 44968 30132
rect 45100 30184 45152 30190
rect 45100 30126 45152 30132
rect 44928 29646 44956 30126
rect 44916 29640 44968 29646
rect 44916 29582 44968 29588
rect 44732 28076 44784 28082
rect 44732 28018 44784 28024
rect 44744 27606 44772 28018
rect 44732 27600 44784 27606
rect 44732 27542 44784 27548
rect 44640 27124 44692 27130
rect 44640 27066 44692 27072
rect 44456 26512 44508 26518
rect 44456 26454 44508 26460
rect 44180 26376 44232 26382
rect 44180 26318 44232 26324
rect 44088 25764 44140 25770
rect 44088 25706 44140 25712
rect 44100 25226 44128 25706
rect 44192 25430 44220 26318
rect 44652 26314 44680 27066
rect 44640 26308 44692 26314
rect 44640 26250 44692 26256
rect 44364 25900 44416 25906
rect 44364 25842 44416 25848
rect 44272 25832 44324 25838
rect 44272 25774 44324 25780
rect 44180 25424 44232 25430
rect 44180 25366 44232 25372
rect 44088 25220 44140 25226
rect 44088 25162 44140 25168
rect 44284 25158 44312 25774
rect 44376 25498 44404 25842
rect 44364 25492 44416 25498
rect 44364 25434 44416 25440
rect 43996 25152 44048 25158
rect 43996 25094 44048 25100
rect 44272 25152 44324 25158
rect 44272 25094 44324 25100
rect 44008 24682 44036 25094
rect 43996 24676 44048 24682
rect 43996 24618 44048 24624
rect 44284 23866 44312 25094
rect 44652 24886 44680 26250
rect 44640 24880 44692 24886
rect 44640 24822 44692 24828
rect 44548 24744 44600 24750
rect 44548 24686 44600 24692
rect 44560 24410 44588 24686
rect 44732 24676 44784 24682
rect 44732 24618 44784 24624
rect 44548 24404 44600 24410
rect 44548 24346 44600 24352
rect 44364 24064 44416 24070
rect 44364 24006 44416 24012
rect 44272 23860 44324 23866
rect 44272 23802 44324 23808
rect 44376 23730 44404 24006
rect 44744 23730 44772 24618
rect 44928 24614 44956 29582
rect 45008 28552 45060 28558
rect 45008 28494 45060 28500
rect 45020 27826 45048 28494
rect 45112 28218 45140 30126
rect 45204 29850 45232 30194
rect 45192 29844 45244 29850
rect 45192 29786 45244 29792
rect 45652 29028 45704 29034
rect 45652 28970 45704 28976
rect 45560 28552 45612 28558
rect 45560 28494 45612 28500
rect 45284 28484 45336 28490
rect 45284 28426 45336 28432
rect 45376 28484 45428 28490
rect 45376 28426 45428 28432
rect 45192 28416 45244 28422
rect 45192 28358 45244 28364
rect 45100 28212 45152 28218
rect 45100 28154 45152 28160
rect 45204 27946 45232 28358
rect 45192 27940 45244 27946
rect 45192 27882 45244 27888
rect 45296 27878 45324 28426
rect 45388 28150 45416 28426
rect 45572 28218 45600 28494
rect 45664 28422 45692 28970
rect 45928 28960 45980 28966
rect 45928 28902 45980 28908
rect 46020 28960 46072 28966
rect 46020 28902 46072 28908
rect 45836 28620 45888 28626
rect 45836 28562 45888 28568
rect 45848 28422 45876 28562
rect 45652 28416 45704 28422
rect 45652 28358 45704 28364
rect 45836 28416 45888 28422
rect 45836 28358 45888 28364
rect 45560 28212 45612 28218
rect 45560 28154 45612 28160
rect 45376 28144 45428 28150
rect 45376 28086 45428 28092
rect 45848 28014 45876 28358
rect 45836 28008 45888 28014
rect 45836 27950 45888 27956
rect 45284 27872 45336 27878
rect 45020 27798 45232 27826
rect 45284 27814 45336 27820
rect 45204 27674 45232 27798
rect 45192 27668 45244 27674
rect 45192 27610 45244 27616
rect 45204 27470 45232 27610
rect 45192 27464 45244 27470
rect 45192 27406 45244 27412
rect 45296 27316 45324 27814
rect 45744 27464 45796 27470
rect 45848 27452 45876 27950
rect 45940 27674 45968 28902
rect 46032 28490 46060 28902
rect 46020 28484 46072 28490
rect 46020 28426 46072 28432
rect 46124 28218 46152 31282
rect 46308 30938 46336 34138
rect 46400 33096 46428 35022
rect 46480 33992 46532 33998
rect 46480 33934 46532 33940
rect 46492 33658 46520 33934
rect 46480 33652 46532 33658
rect 46480 33594 46532 33600
rect 46768 33114 46796 36722
rect 46952 36650 46980 38286
rect 46940 36644 46992 36650
rect 46940 36586 46992 36592
rect 46940 36100 46992 36106
rect 46940 36042 46992 36048
rect 46952 34542 46980 36042
rect 46940 34536 46992 34542
rect 46940 34478 46992 34484
rect 46952 34406 46980 34478
rect 46940 34400 46992 34406
rect 46940 34342 46992 34348
rect 46940 34060 46992 34066
rect 46940 34002 46992 34008
rect 46952 33862 46980 34002
rect 46940 33856 46992 33862
rect 46940 33798 46992 33804
rect 46480 33108 46532 33114
rect 46400 33068 46480 33096
rect 46480 33050 46532 33056
rect 46756 33108 46808 33114
rect 46756 33050 46808 33056
rect 46388 32904 46440 32910
rect 46388 32846 46440 32852
rect 46296 30932 46348 30938
rect 46296 30874 46348 30880
rect 46400 29850 46428 32846
rect 46492 31482 46520 33050
rect 46952 32026 46980 33798
rect 47044 33522 47072 44814
rect 47124 44260 47176 44266
rect 47124 44202 47176 44208
rect 47136 42702 47164 44202
rect 47228 43450 47256 45290
rect 47308 44464 47360 44470
rect 47308 44406 47360 44412
rect 47216 43444 47268 43450
rect 47216 43386 47268 43392
rect 47216 43240 47268 43246
rect 47216 43182 47268 43188
rect 47124 42696 47176 42702
rect 47124 42638 47176 42644
rect 47136 42362 47164 42638
rect 47124 42356 47176 42362
rect 47124 42298 47176 42304
rect 47124 41200 47176 41206
rect 47124 41142 47176 41148
rect 47136 40118 47164 41142
rect 47228 41070 47256 43182
rect 47320 43178 47348 44406
rect 47412 43194 47440 48078
rect 47676 48068 47728 48074
rect 47676 48010 47728 48016
rect 47688 47054 47716 48010
rect 47768 48000 47820 48006
rect 47768 47942 47820 47948
rect 48780 48000 48832 48006
rect 48780 47942 48832 47948
rect 47780 47598 47808 47942
rect 47860 47660 47912 47666
rect 47860 47602 47912 47608
rect 48228 47660 48280 47666
rect 48228 47602 48280 47608
rect 48412 47660 48464 47666
rect 48412 47602 48464 47608
rect 47768 47592 47820 47598
rect 47872 47569 47900 47602
rect 47768 47534 47820 47540
rect 47858 47560 47914 47569
rect 47858 47495 47914 47504
rect 48240 47258 48268 47602
rect 47952 47252 48004 47258
rect 47952 47194 48004 47200
rect 48228 47252 48280 47258
rect 48228 47194 48280 47200
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47860 47048 47912 47054
rect 47860 46990 47912 46996
rect 47768 46980 47820 46986
rect 47768 46922 47820 46928
rect 47780 46510 47808 46922
rect 47676 46504 47728 46510
rect 47676 46446 47728 46452
rect 47768 46504 47820 46510
rect 47768 46446 47820 46452
rect 47584 45892 47636 45898
rect 47584 45834 47636 45840
rect 47596 45286 47624 45834
rect 47688 45422 47716 46446
rect 47780 46170 47808 46446
rect 47768 46164 47820 46170
rect 47768 46106 47820 46112
rect 47768 45484 47820 45490
rect 47768 45426 47820 45432
rect 47676 45416 47728 45422
rect 47676 45358 47728 45364
rect 47492 45280 47544 45286
rect 47492 45222 47544 45228
rect 47584 45280 47636 45286
rect 47584 45222 47636 45228
rect 47504 43314 47532 45222
rect 47688 45082 47716 45358
rect 47676 45076 47728 45082
rect 47676 45018 47728 45024
rect 47676 44192 47728 44198
rect 47676 44134 47728 44140
rect 47582 44024 47638 44033
rect 47582 43959 47638 43968
rect 47596 43790 47624 43959
rect 47584 43784 47636 43790
rect 47584 43726 47636 43732
rect 47688 43314 47716 44134
rect 47780 43897 47808 45426
rect 47872 44538 47900 46990
rect 47964 46170 47992 47194
rect 48320 46980 48372 46986
rect 48320 46922 48372 46928
rect 47952 46164 48004 46170
rect 47952 46106 48004 46112
rect 47952 45824 48004 45830
rect 47952 45766 48004 45772
rect 47860 44532 47912 44538
rect 47860 44474 47912 44480
rect 47766 43888 47822 43897
rect 47766 43823 47822 43832
rect 47492 43308 47544 43314
rect 47492 43250 47544 43256
rect 47676 43308 47728 43314
rect 47676 43250 47728 43256
rect 47308 43172 47360 43178
rect 47412 43166 47532 43194
rect 47308 43114 47360 43120
rect 47320 42702 47348 43114
rect 47308 42696 47360 42702
rect 47308 42638 47360 42644
rect 47308 42084 47360 42090
rect 47308 42026 47360 42032
rect 47320 41546 47348 42026
rect 47308 41540 47360 41546
rect 47308 41482 47360 41488
rect 47400 41472 47452 41478
rect 47400 41414 47452 41420
rect 47412 41138 47440 41414
rect 47400 41132 47452 41138
rect 47400 41074 47452 41080
rect 47216 41064 47268 41070
rect 47216 41006 47268 41012
rect 47124 40112 47176 40118
rect 47124 40054 47176 40060
rect 47136 38010 47164 40054
rect 47228 39642 47256 41006
rect 47400 40928 47452 40934
rect 47400 40870 47452 40876
rect 47412 40526 47440 40870
rect 47400 40520 47452 40526
rect 47400 40462 47452 40468
rect 47504 40458 47532 43166
rect 47780 42344 47808 43823
rect 47860 43648 47912 43654
rect 47860 43590 47912 43596
rect 47872 43246 47900 43590
rect 47860 43240 47912 43246
rect 47860 43182 47912 43188
rect 47780 42316 47900 42344
rect 47768 42220 47820 42226
rect 47768 42162 47820 42168
rect 47676 41676 47728 41682
rect 47780 41664 47808 42162
rect 47872 42090 47900 42316
rect 47860 42084 47912 42090
rect 47860 42026 47912 42032
rect 47964 41750 47992 45766
rect 48134 45520 48190 45529
rect 48134 45455 48190 45464
rect 48228 45484 48280 45490
rect 48148 45422 48176 45455
rect 48228 45426 48280 45432
rect 48136 45416 48188 45422
rect 48136 45358 48188 45364
rect 48240 45354 48268 45426
rect 48228 45348 48280 45354
rect 48228 45290 48280 45296
rect 48240 45082 48268 45290
rect 48228 45076 48280 45082
rect 48228 45018 48280 45024
rect 48228 44872 48280 44878
rect 48228 44814 48280 44820
rect 48240 44538 48268 44814
rect 48228 44532 48280 44538
rect 48228 44474 48280 44480
rect 48332 44402 48360 46922
rect 48424 46374 48452 47602
rect 48792 47598 48820 47942
rect 50294 47900 50602 47920
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47824 50602 47844
rect 48780 47592 48832 47598
rect 48780 47534 48832 47540
rect 48780 47456 48832 47462
rect 48780 47398 48832 47404
rect 48872 47456 48924 47462
rect 48872 47398 48924 47404
rect 48688 46912 48740 46918
rect 48688 46854 48740 46860
rect 48700 46646 48728 46854
rect 48688 46640 48740 46646
rect 48688 46582 48740 46588
rect 48412 46368 48464 46374
rect 48412 46310 48464 46316
rect 48320 44396 48372 44402
rect 48320 44338 48372 44344
rect 48228 44328 48280 44334
rect 48228 44270 48280 44276
rect 48136 43784 48188 43790
rect 48136 43726 48188 43732
rect 48148 43178 48176 43726
rect 48136 43172 48188 43178
rect 48136 43114 48188 43120
rect 48136 42696 48188 42702
rect 48136 42638 48188 42644
rect 47952 41744 48004 41750
rect 47952 41686 48004 41692
rect 47728 41636 47808 41664
rect 47676 41618 47728 41624
rect 47584 40656 47636 40662
rect 47584 40598 47636 40604
rect 47492 40452 47544 40458
rect 47492 40394 47544 40400
rect 47504 39846 47532 40394
rect 47492 39840 47544 39846
rect 47492 39782 47544 39788
rect 47216 39636 47268 39642
rect 47216 39578 47268 39584
rect 47228 39302 47256 39578
rect 47216 39296 47268 39302
rect 47216 39238 47268 39244
rect 47492 38276 47544 38282
rect 47492 38218 47544 38224
rect 47124 38004 47176 38010
rect 47124 37946 47176 37952
rect 47216 37868 47268 37874
rect 47216 37810 47268 37816
rect 47228 37330 47256 37810
rect 47400 37732 47452 37738
rect 47400 37674 47452 37680
rect 47412 37466 47440 37674
rect 47400 37460 47452 37466
rect 47400 37402 47452 37408
rect 47216 37324 47268 37330
rect 47216 37266 47268 37272
rect 47228 35290 47256 37266
rect 47504 37262 47532 38218
rect 47492 37256 47544 37262
rect 47492 37198 47544 37204
rect 47492 36712 47544 36718
rect 47596 36666 47624 40598
rect 47676 40452 47728 40458
rect 47676 40394 47728 40400
rect 47688 40186 47716 40394
rect 47676 40180 47728 40186
rect 47676 40122 47728 40128
rect 47674 37904 47730 37913
rect 47674 37839 47676 37848
rect 47728 37839 47730 37848
rect 47676 37810 47728 37816
rect 47676 37120 47728 37126
rect 47676 37062 47728 37068
rect 47544 36660 47624 36666
rect 47492 36654 47624 36660
rect 47504 36638 47624 36654
rect 47492 36032 47544 36038
rect 47492 35974 47544 35980
rect 47216 35284 47268 35290
rect 47216 35226 47268 35232
rect 47216 35080 47268 35086
rect 47216 35022 47268 35028
rect 47124 34604 47176 34610
rect 47124 34546 47176 34552
rect 47032 33516 47084 33522
rect 47032 33458 47084 33464
rect 47136 33454 47164 34546
rect 47228 34066 47256 35022
rect 47400 35012 47452 35018
rect 47400 34954 47452 34960
rect 47308 34536 47360 34542
rect 47308 34478 47360 34484
rect 47216 34060 47268 34066
rect 47216 34002 47268 34008
rect 47320 33930 47348 34478
rect 47412 33998 47440 34954
rect 47504 34678 47532 35974
rect 47492 34672 47544 34678
rect 47492 34614 47544 34620
rect 47504 34202 47532 34614
rect 47596 34490 47624 36638
rect 47688 36106 47716 37062
rect 47676 36100 47728 36106
rect 47676 36042 47728 36048
rect 47688 34610 47716 36042
rect 47676 34604 47728 34610
rect 47676 34546 47728 34552
rect 47596 34462 47716 34490
rect 47492 34196 47544 34202
rect 47492 34138 47544 34144
rect 47584 34196 47636 34202
rect 47584 34138 47636 34144
rect 47400 33992 47452 33998
rect 47400 33934 47452 33940
rect 47308 33924 47360 33930
rect 47308 33866 47360 33872
rect 47216 33856 47268 33862
rect 47216 33798 47268 33804
rect 47228 33658 47256 33798
rect 47320 33658 47348 33866
rect 47216 33652 47268 33658
rect 47216 33594 47268 33600
rect 47308 33652 47360 33658
rect 47308 33594 47360 33600
rect 47124 33448 47176 33454
rect 47124 33390 47176 33396
rect 47136 33114 47164 33390
rect 47124 33108 47176 33114
rect 47124 33050 47176 33056
rect 46940 32020 46992 32026
rect 46940 31962 46992 31968
rect 46756 31952 46808 31958
rect 46756 31894 46808 31900
rect 46664 31884 46716 31890
rect 46664 31826 46716 31832
rect 46676 31754 46704 31826
rect 46768 31822 46796 31894
rect 46756 31816 46808 31822
rect 46756 31758 46808 31764
rect 46584 31726 46704 31754
rect 46480 31476 46532 31482
rect 46480 31418 46532 31424
rect 46480 30728 46532 30734
rect 46480 30670 46532 30676
rect 46388 29844 46440 29850
rect 46388 29786 46440 29792
rect 46492 29102 46520 30670
rect 46584 30598 46612 31726
rect 46768 30734 46796 31758
rect 47124 31680 47176 31686
rect 47124 31622 47176 31628
rect 47136 30734 47164 31622
rect 46756 30728 46808 30734
rect 46756 30670 46808 30676
rect 47124 30728 47176 30734
rect 47124 30670 47176 30676
rect 46572 30592 46624 30598
rect 46572 30534 46624 30540
rect 46584 29578 46612 30534
rect 46768 30258 46796 30670
rect 46756 30252 46808 30258
rect 46756 30194 46808 30200
rect 46768 29782 46796 30194
rect 46756 29776 46808 29782
rect 46756 29718 46808 29724
rect 46572 29572 46624 29578
rect 46572 29514 46624 29520
rect 46664 29164 46716 29170
rect 46664 29106 46716 29112
rect 46480 29096 46532 29102
rect 46480 29038 46532 29044
rect 46112 28212 46164 28218
rect 46112 28154 46164 28160
rect 46492 28082 46520 29038
rect 46676 28082 46704 29106
rect 47228 28558 47256 33594
rect 47308 33516 47360 33522
rect 47308 33458 47360 33464
rect 47320 31686 47348 33458
rect 47412 32570 47440 33934
rect 47504 33522 47532 34138
rect 47492 33516 47544 33522
rect 47492 33458 47544 33464
rect 47596 33318 47624 34138
rect 47584 33312 47636 33318
rect 47584 33254 47636 33260
rect 47492 32904 47544 32910
rect 47492 32846 47544 32852
rect 47400 32564 47452 32570
rect 47400 32506 47452 32512
rect 47308 31680 47360 31686
rect 47308 31622 47360 31628
rect 47504 28762 47532 32846
rect 47584 31340 47636 31346
rect 47584 31282 47636 31288
rect 47596 29850 47624 31282
rect 47584 29844 47636 29850
rect 47584 29786 47636 29792
rect 47584 29640 47636 29646
rect 47584 29582 47636 29588
rect 47492 28756 47544 28762
rect 47492 28698 47544 28704
rect 47216 28552 47268 28558
rect 47216 28494 47268 28500
rect 47228 28150 47256 28494
rect 47216 28144 47268 28150
rect 47216 28086 47268 28092
rect 46388 28076 46440 28082
rect 46388 28018 46440 28024
rect 46480 28076 46532 28082
rect 46480 28018 46532 28024
rect 46664 28076 46716 28082
rect 46664 28018 46716 28024
rect 46400 27674 46428 28018
rect 45928 27668 45980 27674
rect 45928 27610 45980 27616
rect 46388 27668 46440 27674
rect 46388 27610 46440 27616
rect 45796 27424 45876 27452
rect 45928 27464 45980 27470
rect 45744 27406 45796 27412
rect 45928 27406 45980 27412
rect 46296 27464 46348 27470
rect 46296 27406 46348 27412
rect 45940 27334 45968 27406
rect 45376 27328 45428 27334
rect 45296 27288 45376 27316
rect 45376 27270 45428 27276
rect 45928 27328 45980 27334
rect 45928 27270 45980 27276
rect 46308 26994 46336 27406
rect 46296 26988 46348 26994
rect 46296 26930 46348 26936
rect 46308 26042 46336 26930
rect 46388 26308 46440 26314
rect 46388 26250 46440 26256
rect 46296 26036 46348 26042
rect 46296 25978 46348 25984
rect 45284 25492 45336 25498
rect 45284 25434 45336 25440
rect 45192 25152 45244 25158
rect 45192 25094 45244 25100
rect 45204 24954 45232 25094
rect 45192 24948 45244 24954
rect 45192 24890 45244 24896
rect 45296 24818 45324 25434
rect 46296 24880 46348 24886
rect 46400 24857 46428 26250
rect 46296 24822 46348 24828
rect 46386 24848 46442 24857
rect 45284 24812 45336 24818
rect 45284 24754 45336 24760
rect 45468 24676 45520 24682
rect 45468 24618 45520 24624
rect 44916 24608 44968 24614
rect 44916 24550 44968 24556
rect 45192 24200 45244 24206
rect 45192 24142 45244 24148
rect 45204 23866 45232 24142
rect 45480 24070 45508 24618
rect 45744 24608 45796 24614
rect 45744 24550 45796 24556
rect 45836 24608 45888 24614
rect 45836 24550 45888 24556
rect 45756 24274 45784 24550
rect 45848 24342 45876 24550
rect 45836 24336 45888 24342
rect 45836 24278 45888 24284
rect 46308 24274 46336 24822
rect 46386 24783 46388 24792
rect 46440 24783 46442 24792
rect 46388 24754 46440 24760
rect 45744 24268 45796 24274
rect 45744 24210 45796 24216
rect 46296 24268 46348 24274
rect 46296 24210 46348 24216
rect 45928 24200 45980 24206
rect 45928 24142 45980 24148
rect 45468 24064 45520 24070
rect 45468 24006 45520 24012
rect 45480 23866 45508 24006
rect 45192 23860 45244 23866
rect 45192 23802 45244 23808
rect 45468 23860 45520 23866
rect 45468 23802 45520 23808
rect 45480 23730 45508 23802
rect 45940 23730 45968 24142
rect 44364 23724 44416 23730
rect 44364 23666 44416 23672
rect 44640 23724 44692 23730
rect 44640 23666 44692 23672
rect 44732 23724 44784 23730
rect 44732 23666 44784 23672
rect 45468 23724 45520 23730
rect 45468 23666 45520 23672
rect 45928 23724 45980 23730
rect 45928 23666 45980 23672
rect 44272 23588 44324 23594
rect 44272 23530 44324 23536
rect 43904 23316 43956 23322
rect 43904 23258 43956 23264
rect 44284 23118 44312 23530
rect 44376 23186 44404 23666
rect 44652 23526 44680 23666
rect 45652 23656 45704 23662
rect 45652 23598 45704 23604
rect 45664 23526 45692 23598
rect 44640 23520 44692 23526
rect 44640 23462 44692 23468
rect 45652 23520 45704 23526
rect 45652 23462 45704 23468
rect 44364 23180 44416 23186
rect 44364 23122 44416 23128
rect 44272 23112 44324 23118
rect 44272 23054 44324 23060
rect 44364 22976 44416 22982
rect 44364 22918 44416 22924
rect 44376 22642 44404 22918
rect 44364 22636 44416 22642
rect 44364 22578 44416 22584
rect 44272 22500 44324 22506
rect 44272 22442 44324 22448
rect 43812 22092 43864 22098
rect 43812 22034 43864 22040
rect 43824 21962 43852 22034
rect 43536 21956 43588 21962
rect 43536 21898 43588 21904
rect 43812 21956 43864 21962
rect 43812 21898 43864 21904
rect 44284 21894 44312 22442
rect 44652 22234 44680 23462
rect 46308 23186 46336 24210
rect 46400 23798 46428 24754
rect 46492 24410 46520 28018
rect 47124 26920 47176 26926
rect 47124 26862 47176 26868
rect 47136 26586 47164 26862
rect 47228 26586 47256 28086
rect 47504 28014 47532 28698
rect 47596 28422 47624 29582
rect 47584 28416 47636 28422
rect 47584 28358 47636 28364
rect 47492 28008 47544 28014
rect 47492 27950 47544 27956
rect 47688 27538 47716 34462
rect 47780 30666 47808 41636
rect 47964 40730 47992 41686
rect 47952 40724 48004 40730
rect 47952 40666 48004 40672
rect 47860 40656 47912 40662
rect 47860 40598 47912 40604
rect 47872 40526 47900 40598
rect 47860 40520 47912 40526
rect 47860 40462 47912 40468
rect 47952 40520 48004 40526
rect 47952 40462 48004 40468
rect 47860 37664 47912 37670
rect 47860 37606 47912 37612
rect 47872 37466 47900 37606
rect 47860 37460 47912 37466
rect 47860 37402 47912 37408
rect 47964 34490 47992 40462
rect 48148 40458 48176 42638
rect 48240 42566 48268 44270
rect 48320 42696 48372 42702
rect 48320 42638 48372 42644
rect 48228 42560 48280 42566
rect 48228 42502 48280 42508
rect 48240 41138 48268 42502
rect 48332 41818 48360 42638
rect 48320 41812 48372 41818
rect 48320 41754 48372 41760
rect 48424 41698 48452 46310
rect 48792 45558 48820 47398
rect 48884 47054 48912 47398
rect 48872 47048 48924 47054
rect 48872 46990 48924 46996
rect 49884 47048 49936 47054
rect 49884 46990 49936 46996
rect 49976 47048 50028 47054
rect 49976 46990 50028 46996
rect 49792 46980 49844 46986
rect 49792 46922 49844 46928
rect 49608 46912 49660 46918
rect 49608 46854 49660 46860
rect 49620 45558 49648 46854
rect 49804 46578 49832 46922
rect 49792 46572 49844 46578
rect 49792 46514 49844 46520
rect 48780 45552 48832 45558
rect 48780 45494 48832 45500
rect 49608 45552 49660 45558
rect 49608 45494 49660 45500
rect 48964 45484 49016 45490
rect 48964 45426 49016 45432
rect 48976 44538 49004 45426
rect 49056 45348 49108 45354
rect 49056 45290 49108 45296
rect 49068 44946 49096 45290
rect 49516 45076 49568 45082
rect 49516 45018 49568 45024
rect 49424 45008 49476 45014
rect 49422 44976 49424 44985
rect 49476 44976 49478 44985
rect 49056 44940 49108 44946
rect 49056 44882 49108 44888
rect 49332 44940 49384 44946
rect 49528 44946 49556 45018
rect 49422 44911 49478 44920
rect 49516 44940 49568 44946
rect 49332 44882 49384 44888
rect 49516 44882 49568 44888
rect 48964 44532 49016 44538
rect 48964 44474 49016 44480
rect 49344 44402 49372 44882
rect 49424 44872 49476 44878
rect 49424 44814 49476 44820
rect 49436 44470 49464 44814
rect 49424 44464 49476 44470
rect 49424 44406 49476 44412
rect 48780 44396 48832 44402
rect 48780 44338 48832 44344
rect 49332 44396 49384 44402
rect 49332 44338 49384 44344
rect 48596 43784 48648 43790
rect 48596 43726 48648 43732
rect 48608 42294 48636 43726
rect 48596 42288 48648 42294
rect 48596 42230 48648 42236
rect 48504 42220 48556 42226
rect 48504 42162 48556 42168
rect 48332 41670 48452 41698
rect 48228 41132 48280 41138
rect 48228 41074 48280 41080
rect 48136 40452 48188 40458
rect 48136 40394 48188 40400
rect 48240 40338 48268 41074
rect 48332 40576 48360 41670
rect 48516 41614 48544 42162
rect 48504 41608 48556 41614
rect 48504 41550 48556 41556
rect 48688 41064 48740 41070
rect 48688 41006 48740 41012
rect 48412 40588 48464 40594
rect 48332 40548 48412 40576
rect 48412 40530 48464 40536
rect 48056 40310 48268 40338
rect 48056 38962 48084 40310
rect 48318 39944 48374 39953
rect 48318 39879 48320 39888
rect 48372 39879 48374 39888
rect 48320 39850 48372 39856
rect 48700 39438 48728 41006
rect 48792 40118 48820 44338
rect 49344 43926 49372 44338
rect 49332 43920 49384 43926
rect 49332 43862 49384 43868
rect 49620 43858 49648 45494
rect 49700 45484 49752 45490
rect 49700 45426 49752 45432
rect 49712 45082 49740 45426
rect 49700 45076 49752 45082
rect 49700 45018 49752 45024
rect 49700 44736 49752 44742
rect 49700 44678 49752 44684
rect 49712 44441 49740 44678
rect 49698 44432 49754 44441
rect 49698 44367 49754 44376
rect 49608 43852 49660 43858
rect 49608 43794 49660 43800
rect 49804 42906 49832 46514
rect 49896 46374 49924 46990
rect 49988 46918 50016 46990
rect 49976 46912 50028 46918
rect 49976 46854 50028 46860
rect 50068 46912 50120 46918
rect 50068 46854 50120 46860
rect 50080 46714 50108 46854
rect 50294 46812 50602 46832
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46736 50602 46756
rect 50068 46708 50120 46714
rect 50068 46650 50120 46656
rect 50080 46578 50108 46650
rect 50068 46572 50120 46578
rect 50068 46514 50120 46520
rect 50712 46572 50764 46578
rect 50712 46514 50764 46520
rect 49884 46368 49936 46374
rect 49884 46310 49936 46316
rect 49884 46096 49936 46102
rect 49884 46038 49936 46044
rect 49792 42900 49844 42906
rect 49792 42842 49844 42848
rect 49240 42356 49292 42362
rect 49240 42298 49292 42304
rect 48872 42220 48924 42226
rect 48872 42162 48924 42168
rect 48884 40186 48912 42162
rect 49252 41274 49280 42298
rect 49792 42152 49844 42158
rect 49792 42094 49844 42100
rect 49240 41268 49292 41274
rect 49240 41210 49292 41216
rect 49608 41200 49660 41206
rect 49608 41142 49660 41148
rect 49240 41132 49292 41138
rect 49240 41074 49292 41080
rect 48872 40180 48924 40186
rect 48872 40122 48924 40128
rect 48780 40112 48832 40118
rect 48780 40054 48832 40060
rect 48596 39432 48648 39438
rect 48596 39374 48648 39380
rect 48688 39432 48740 39438
rect 48688 39374 48740 39380
rect 48504 39024 48556 39030
rect 48504 38966 48556 38972
rect 48044 38956 48096 38962
rect 48044 38898 48096 38904
rect 48056 37074 48084 38898
rect 48412 38888 48464 38894
rect 48412 38830 48464 38836
rect 48424 38350 48452 38830
rect 48412 38344 48464 38350
rect 48412 38286 48464 38292
rect 48320 38208 48372 38214
rect 48320 38150 48372 38156
rect 48136 37664 48188 37670
rect 48136 37606 48188 37612
rect 48148 37398 48176 37606
rect 48136 37392 48188 37398
rect 48136 37334 48188 37340
rect 48148 37262 48176 37334
rect 48136 37256 48188 37262
rect 48136 37198 48188 37204
rect 48332 37194 48360 38150
rect 48516 37262 48544 38966
rect 48608 38196 48636 39374
rect 48700 38758 48728 39374
rect 48792 39030 48820 40054
rect 48780 39024 48832 39030
rect 48780 38966 48832 38972
rect 48688 38752 48740 38758
rect 48688 38694 48740 38700
rect 48884 38350 48912 40122
rect 49252 40118 49280 41074
rect 49516 40996 49568 41002
rect 49516 40938 49568 40944
rect 49424 40928 49476 40934
rect 49424 40870 49476 40876
rect 49332 40520 49384 40526
rect 49332 40462 49384 40468
rect 49240 40112 49292 40118
rect 49240 40054 49292 40060
rect 48964 39432 49016 39438
rect 48964 39374 49016 39380
rect 48976 38894 49004 39374
rect 49252 39098 49280 40054
rect 49344 39846 49372 40462
rect 49332 39840 49384 39846
rect 49332 39782 49384 39788
rect 49344 39574 49372 39782
rect 49332 39568 49384 39574
rect 49332 39510 49384 39516
rect 49240 39092 49292 39098
rect 49240 39034 49292 39040
rect 48964 38888 49016 38894
rect 48964 38830 49016 38836
rect 48964 38752 49016 38758
rect 48964 38694 49016 38700
rect 48872 38344 48924 38350
rect 48872 38286 48924 38292
rect 48608 38168 48728 38196
rect 48596 37868 48648 37874
rect 48596 37810 48648 37816
rect 48504 37256 48556 37262
rect 48504 37198 48556 37204
rect 48320 37188 48372 37194
rect 48320 37130 48372 37136
rect 48412 37188 48464 37194
rect 48412 37130 48464 37136
rect 48136 37120 48188 37126
rect 48056 37068 48136 37074
rect 48056 37062 48188 37068
rect 48056 37046 48176 37062
rect 48148 36718 48176 37046
rect 48136 36712 48188 36718
rect 48136 36654 48188 36660
rect 48044 36576 48096 36582
rect 48044 36518 48096 36524
rect 48056 36242 48084 36518
rect 48044 36236 48096 36242
rect 48044 36178 48096 36184
rect 48228 36168 48280 36174
rect 48228 36110 48280 36116
rect 47872 34462 47992 34490
rect 47872 33998 47900 34462
rect 48240 34406 48268 36110
rect 47952 34400 48004 34406
rect 47952 34342 48004 34348
rect 48228 34400 48280 34406
rect 48228 34342 48280 34348
rect 47860 33992 47912 33998
rect 47860 33934 47912 33940
rect 47964 33522 47992 34342
rect 48332 34066 48360 37130
rect 48424 35698 48452 37130
rect 48608 36854 48636 37810
rect 48596 36848 48648 36854
rect 48596 36790 48648 36796
rect 48608 35834 48636 36790
rect 48596 35828 48648 35834
rect 48596 35770 48648 35776
rect 48700 35714 48728 38168
rect 48884 37738 48912 38286
rect 48872 37732 48924 37738
rect 48872 37674 48924 37680
rect 48780 36780 48832 36786
rect 48780 36722 48832 36728
rect 48412 35692 48464 35698
rect 48412 35634 48464 35640
rect 48516 35686 48728 35714
rect 48412 34604 48464 34610
rect 48412 34546 48464 34552
rect 48320 34060 48372 34066
rect 48320 34002 48372 34008
rect 48424 33998 48452 34546
rect 48412 33992 48464 33998
rect 48412 33934 48464 33940
rect 48412 33856 48464 33862
rect 48412 33798 48464 33804
rect 48424 33658 48452 33798
rect 48412 33652 48464 33658
rect 48412 33594 48464 33600
rect 47952 33516 48004 33522
rect 47952 33458 48004 33464
rect 47964 33046 47992 33458
rect 48424 33266 48452 33594
rect 48056 33238 48452 33266
rect 48056 33114 48084 33238
rect 48044 33108 48096 33114
rect 48044 33050 48096 33056
rect 48136 33108 48188 33114
rect 48136 33050 48188 33056
rect 47952 33040 48004 33046
rect 47952 32982 48004 32988
rect 47860 32972 47912 32978
rect 47860 32914 47912 32920
rect 47872 32298 47900 32914
rect 47952 32768 48004 32774
rect 48148 32756 48176 33050
rect 48004 32728 48176 32756
rect 47952 32710 48004 32716
rect 48044 32428 48096 32434
rect 48044 32370 48096 32376
rect 47860 32292 47912 32298
rect 47860 32234 47912 32240
rect 47952 31816 48004 31822
rect 47952 31758 48004 31764
rect 47964 30938 47992 31758
rect 48056 31346 48084 32370
rect 48148 31482 48176 32728
rect 48320 32564 48372 32570
rect 48320 32506 48372 32512
rect 48228 32428 48280 32434
rect 48228 32370 48280 32376
rect 48136 31476 48188 31482
rect 48136 31418 48188 31424
rect 48044 31340 48096 31346
rect 48044 31282 48096 31288
rect 48240 31142 48268 32370
rect 48332 31958 48360 32506
rect 48320 31952 48372 31958
rect 48320 31894 48372 31900
rect 48228 31136 48280 31142
rect 48228 31078 48280 31084
rect 47952 30932 48004 30938
rect 47952 30874 48004 30880
rect 47768 30660 47820 30666
rect 47768 30602 47820 30608
rect 47964 30258 47992 30874
rect 47952 30252 48004 30258
rect 47952 30194 48004 30200
rect 48136 30048 48188 30054
rect 48136 29990 48188 29996
rect 47860 29776 47912 29782
rect 47860 29718 47912 29724
rect 47768 29572 47820 29578
rect 47768 29514 47820 29520
rect 47780 28558 47808 29514
rect 47872 28558 47900 29718
rect 48148 29646 48176 29990
rect 48136 29640 48188 29646
rect 48136 29582 48188 29588
rect 48516 28966 48544 35686
rect 48596 35624 48648 35630
rect 48596 35566 48648 35572
rect 48608 33658 48636 35566
rect 48688 35216 48740 35222
rect 48688 35158 48740 35164
rect 48700 34610 48728 35158
rect 48688 34604 48740 34610
rect 48688 34546 48740 34552
rect 48596 33652 48648 33658
rect 48596 33594 48648 33600
rect 48688 32496 48740 32502
rect 48688 32438 48740 32444
rect 48700 32026 48728 32438
rect 48688 32020 48740 32026
rect 48688 31962 48740 31968
rect 48792 30870 48820 36722
rect 48884 32434 48912 37674
rect 48976 36582 49004 38694
rect 49056 38480 49108 38486
rect 49056 38422 49108 38428
rect 49068 37874 49096 38422
rect 49056 37868 49108 37874
rect 49056 37810 49108 37816
rect 49056 37324 49108 37330
rect 49056 37266 49108 37272
rect 48964 36576 49016 36582
rect 48964 36518 49016 36524
rect 49068 35494 49096 37266
rect 49148 36848 49200 36854
rect 49148 36790 49200 36796
rect 49056 35488 49108 35494
rect 49056 35430 49108 35436
rect 49068 35290 49096 35430
rect 49056 35284 49108 35290
rect 49056 35226 49108 35232
rect 48964 35012 49016 35018
rect 48964 34954 49016 34960
rect 48976 33504 49004 34954
rect 49056 34604 49108 34610
rect 49056 34546 49108 34552
rect 49068 33969 49096 34546
rect 49054 33960 49110 33969
rect 49054 33895 49110 33904
rect 49056 33516 49108 33522
rect 48976 33476 49056 33504
rect 49056 33458 49108 33464
rect 49068 33289 49096 33458
rect 49054 33280 49110 33289
rect 49054 33215 49110 33224
rect 48872 32428 48924 32434
rect 48872 32370 48924 32376
rect 48884 32026 48912 32370
rect 48872 32020 48924 32026
rect 48872 31962 48924 31968
rect 49160 30938 49188 36790
rect 49344 35766 49372 39510
rect 49436 39302 49464 40870
rect 49528 40730 49556 40938
rect 49620 40730 49648 41142
rect 49516 40724 49568 40730
rect 49516 40666 49568 40672
rect 49608 40724 49660 40730
rect 49608 40666 49660 40672
rect 49424 39296 49476 39302
rect 49424 39238 49476 39244
rect 49700 38888 49752 38894
rect 49700 38830 49752 38836
rect 49712 38434 49740 38830
rect 49620 38406 49740 38434
rect 49516 37868 49568 37874
rect 49516 37810 49568 37816
rect 49528 37330 49556 37810
rect 49516 37324 49568 37330
rect 49516 37266 49568 37272
rect 49424 36576 49476 36582
rect 49424 36518 49476 36524
rect 49332 35760 49384 35766
rect 49332 35702 49384 35708
rect 49240 35692 49292 35698
rect 49240 35634 49292 35640
rect 49252 34542 49280 35634
rect 49240 34536 49292 34542
rect 49240 34478 49292 34484
rect 49252 33522 49280 34478
rect 49332 33924 49384 33930
rect 49332 33866 49384 33872
rect 49240 33516 49292 33522
rect 49240 33458 49292 33464
rect 49252 33425 49280 33458
rect 49238 33416 49294 33425
rect 49344 33386 49372 33866
rect 49238 33351 49294 33360
rect 49332 33380 49384 33386
rect 49332 33322 49384 33328
rect 49240 32836 49292 32842
rect 49240 32778 49292 32784
rect 49252 31414 49280 32778
rect 49436 31958 49464 36518
rect 49424 31952 49476 31958
rect 49424 31894 49476 31900
rect 49528 31754 49556 37266
rect 49620 36718 49648 38406
rect 49700 38344 49752 38350
rect 49700 38286 49752 38292
rect 49712 38010 49740 38286
rect 49804 38049 49832 42094
rect 49896 40662 49924 46038
rect 50160 45960 50212 45966
rect 50160 45902 50212 45908
rect 50068 44396 50120 44402
rect 50068 44338 50120 44344
rect 50080 43994 50108 44338
rect 50068 43988 50120 43994
rect 50068 43930 50120 43936
rect 50068 43784 50120 43790
rect 50068 43726 50120 43732
rect 49976 43308 50028 43314
rect 49976 43250 50028 43256
rect 49988 42702 50016 43250
rect 50080 43246 50108 43726
rect 50068 43240 50120 43246
rect 50068 43182 50120 43188
rect 49976 42696 50028 42702
rect 49976 42638 50028 42644
rect 49988 42226 50016 42638
rect 50080 42362 50108 43182
rect 50068 42356 50120 42362
rect 50068 42298 50120 42304
rect 49976 42220 50028 42226
rect 49976 42162 50028 42168
rect 49884 40656 49936 40662
rect 49884 40598 49936 40604
rect 49884 40044 49936 40050
rect 49884 39986 49936 39992
rect 49896 38894 49924 39986
rect 49884 38888 49936 38894
rect 49884 38830 49936 38836
rect 49988 38554 50016 42162
rect 50172 42090 50200 45902
rect 50724 45830 50752 46514
rect 51264 46504 51316 46510
rect 51264 46446 51316 46452
rect 50988 46368 51040 46374
rect 50988 46310 51040 46316
rect 51000 45966 51028 46310
rect 51276 45966 51304 46446
rect 50988 45960 51040 45966
rect 50988 45902 51040 45908
rect 51264 45960 51316 45966
rect 51264 45902 51316 45908
rect 51816 45960 51868 45966
rect 51816 45902 51868 45908
rect 50712 45824 50764 45830
rect 50712 45766 50764 45772
rect 50294 45724 50602 45744
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45648 50602 45668
rect 50724 45082 50752 45766
rect 51448 45484 51500 45490
rect 51448 45426 51500 45432
rect 51356 45416 51408 45422
rect 51356 45358 51408 45364
rect 51368 45082 51396 45358
rect 50712 45076 50764 45082
rect 50712 45018 50764 45024
rect 51356 45076 51408 45082
rect 51356 45018 51408 45024
rect 50896 44736 50948 44742
rect 50896 44678 50948 44684
rect 50294 44636 50602 44656
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44560 50602 44580
rect 50908 44538 50936 44678
rect 50896 44532 50948 44538
rect 50896 44474 50948 44480
rect 51460 44470 51488 45426
rect 51828 45422 51856 45902
rect 52092 45892 52144 45898
rect 52092 45834 52144 45840
rect 51816 45416 51868 45422
rect 51816 45358 51868 45364
rect 52000 45348 52052 45354
rect 52000 45290 52052 45296
rect 50988 44464 51040 44470
rect 50988 44406 51040 44412
rect 51448 44464 51500 44470
rect 51448 44406 51500 44412
rect 50896 44328 50948 44334
rect 50896 44270 50948 44276
rect 50620 43784 50672 43790
rect 50804 43784 50856 43790
rect 50672 43732 50752 43738
rect 50620 43726 50752 43732
rect 50804 43726 50856 43732
rect 50632 43710 50752 43726
rect 50620 43648 50672 43654
rect 50620 43590 50672 43596
rect 50294 43548 50602 43568
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43472 50602 43492
rect 50632 43246 50660 43590
rect 50724 43450 50752 43710
rect 50816 43450 50844 43726
rect 50712 43444 50764 43450
rect 50712 43386 50764 43392
rect 50804 43444 50856 43450
rect 50804 43386 50856 43392
rect 50620 43240 50672 43246
rect 50620 43182 50672 43188
rect 50632 42634 50660 43182
rect 50620 42628 50672 42634
rect 50620 42570 50672 42576
rect 50294 42460 50602 42480
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42384 50602 42404
rect 50160 42084 50212 42090
rect 50160 42026 50212 42032
rect 50068 41608 50120 41614
rect 50068 41550 50120 41556
rect 50080 41138 50108 41550
rect 50294 41372 50602 41392
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41296 50602 41316
rect 50068 41132 50120 41138
rect 50068 41074 50120 41080
rect 50528 41064 50580 41070
rect 50528 41006 50580 41012
rect 50540 40594 50568 41006
rect 50068 40588 50120 40594
rect 50068 40530 50120 40536
rect 50528 40588 50580 40594
rect 50528 40530 50580 40536
rect 50080 39370 50108 40530
rect 50294 40284 50602 40304
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40208 50602 40228
rect 50068 39364 50120 39370
rect 50068 39306 50120 39312
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 50632 38962 50660 42570
rect 50724 41614 50752 43386
rect 50908 43178 50936 44270
rect 51000 43858 51028 44406
rect 52012 44282 52040 45290
rect 52104 44878 52132 45834
rect 52736 45280 52788 45286
rect 52736 45222 52788 45228
rect 52644 44940 52696 44946
rect 52644 44882 52696 44888
rect 52092 44872 52144 44878
rect 52092 44814 52144 44820
rect 52104 44402 52132 44814
rect 52092 44396 52144 44402
rect 52092 44338 52144 44344
rect 52656 44334 52684 44882
rect 52748 44878 52776 45222
rect 55496 45008 55548 45014
rect 55494 44976 55496 44985
rect 55548 44976 55550 44985
rect 53840 44940 53892 44946
rect 55494 44911 55550 44920
rect 53840 44882 53892 44888
rect 52736 44872 52788 44878
rect 52736 44814 52788 44820
rect 53656 44872 53708 44878
rect 53656 44814 53708 44820
rect 52920 44736 52972 44742
rect 52920 44678 52972 44684
rect 52932 44538 52960 44678
rect 53668 44538 53696 44814
rect 52920 44532 52972 44538
rect 52920 44474 52972 44480
rect 53656 44532 53708 44538
rect 53656 44474 53708 44480
rect 53852 44334 53880 44882
rect 55128 44464 55180 44470
rect 55128 44406 55180 44412
rect 52644 44328 52696 44334
rect 52012 44266 52132 44282
rect 52644 44270 52696 44276
rect 53840 44328 53892 44334
rect 53840 44270 53892 44276
rect 52012 44260 52144 44266
rect 52012 44254 52092 44260
rect 52092 44202 52144 44208
rect 50988 43852 51040 43858
rect 50988 43794 51040 43800
rect 51448 43308 51500 43314
rect 51448 43250 51500 43256
rect 50896 43172 50948 43178
rect 50896 43114 50948 43120
rect 51460 42906 51488 43250
rect 51448 42900 51500 42906
rect 51448 42842 51500 42848
rect 50804 42628 50856 42634
rect 50804 42570 50856 42576
rect 50816 42226 50844 42570
rect 51540 42560 51592 42566
rect 51540 42502 51592 42508
rect 51552 42226 51580 42502
rect 50804 42220 50856 42226
rect 50804 42162 50856 42168
rect 51540 42220 51592 42226
rect 51540 42162 51592 42168
rect 51908 42220 51960 42226
rect 51908 42162 51960 42168
rect 50804 42084 50856 42090
rect 50804 42026 50856 42032
rect 50712 41608 50764 41614
rect 50712 41550 50764 41556
rect 50724 38978 50752 41550
rect 50816 40050 50844 42026
rect 51080 41676 51132 41682
rect 51080 41618 51132 41624
rect 51092 41478 51120 41618
rect 51172 41608 51224 41614
rect 51172 41550 51224 41556
rect 50988 41472 51040 41478
rect 50988 41414 51040 41420
rect 51080 41472 51132 41478
rect 51080 41414 51132 41420
rect 51000 41138 51028 41414
rect 51184 41274 51212 41550
rect 51448 41472 51500 41478
rect 51448 41414 51500 41420
rect 51172 41268 51224 41274
rect 51172 41210 51224 41216
rect 50988 41132 51040 41138
rect 50988 41074 51040 41080
rect 51080 40996 51132 41002
rect 51080 40938 51132 40944
rect 51092 40186 51120 40938
rect 51184 40458 51212 41210
rect 51460 40526 51488 41414
rect 51552 41274 51580 42162
rect 51540 41268 51592 41274
rect 51540 41210 51592 41216
rect 51920 41206 51948 42162
rect 51908 41200 51960 41206
rect 51908 41142 51960 41148
rect 51632 40928 51684 40934
rect 51632 40870 51684 40876
rect 51540 40656 51592 40662
rect 51540 40598 51592 40604
rect 51448 40520 51500 40526
rect 51448 40462 51500 40468
rect 51172 40452 51224 40458
rect 51172 40394 51224 40400
rect 51080 40180 51132 40186
rect 51080 40122 51132 40128
rect 51184 40050 51212 40394
rect 51264 40384 51316 40390
rect 51264 40326 51316 40332
rect 50804 40044 50856 40050
rect 50804 39986 50856 39992
rect 51172 40044 51224 40050
rect 51172 39986 51224 39992
rect 50816 39302 50844 39986
rect 51184 39506 51212 39986
rect 51172 39500 51224 39506
rect 51172 39442 51224 39448
rect 50804 39296 50856 39302
rect 50804 39238 50856 39244
rect 51172 39296 51224 39302
rect 51172 39238 51224 39244
rect 50620 38956 50672 38962
rect 50724 38950 50936 38978
rect 50620 38898 50672 38904
rect 49976 38548 50028 38554
rect 49976 38490 50028 38496
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 49790 38040 49846 38049
rect 49700 38004 49752 38010
rect 50294 38032 50602 38052
rect 49790 37975 49846 37984
rect 49700 37946 49752 37952
rect 50632 37874 50660 38898
rect 50712 38888 50764 38894
rect 50712 38830 50764 38836
rect 50724 38282 50752 38830
rect 50712 38276 50764 38282
rect 50712 38218 50764 38224
rect 50724 37942 50752 38218
rect 50712 37936 50764 37942
rect 50712 37878 50764 37884
rect 49792 37868 49844 37874
rect 49792 37810 49844 37816
rect 49976 37868 50028 37874
rect 49976 37810 50028 37816
rect 50068 37868 50120 37874
rect 50068 37810 50120 37816
rect 50252 37868 50304 37874
rect 50252 37810 50304 37816
rect 50620 37868 50672 37874
rect 50620 37810 50672 37816
rect 49700 37324 49752 37330
rect 49700 37266 49752 37272
rect 49608 36712 49660 36718
rect 49608 36654 49660 36660
rect 49620 32774 49648 36654
rect 49608 32768 49660 32774
rect 49608 32710 49660 32716
rect 49344 31726 49556 31754
rect 49240 31408 49292 31414
rect 49240 31350 49292 31356
rect 49344 31346 49372 31726
rect 49712 31482 49740 37266
rect 49804 36854 49832 37810
rect 49884 37800 49936 37806
rect 49884 37742 49936 37748
rect 49792 36848 49844 36854
rect 49792 36790 49844 36796
rect 49896 36666 49924 37742
rect 49988 37126 50016 37810
rect 49976 37120 50028 37126
rect 49976 37062 50028 37068
rect 49804 36638 49924 36666
rect 49804 31754 49832 36638
rect 49988 36582 50016 37062
rect 50080 36854 50108 37810
rect 50160 37664 50212 37670
rect 50160 37606 50212 37612
rect 50068 36848 50120 36854
rect 50068 36790 50120 36796
rect 50172 36786 50200 37606
rect 50264 37262 50292 37810
rect 50620 37732 50672 37738
rect 50620 37674 50672 37680
rect 50632 37262 50660 37674
rect 50252 37256 50304 37262
rect 50252 37198 50304 37204
rect 50620 37256 50672 37262
rect 50620 37198 50672 37204
rect 50724 37074 50752 37878
rect 50632 37046 50752 37074
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50160 36780 50212 36786
rect 50160 36722 50212 36728
rect 49976 36576 50028 36582
rect 49976 36518 50028 36524
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 49884 35760 49936 35766
rect 49884 35702 49936 35708
rect 49896 35057 49924 35702
rect 50632 35494 50660 37046
rect 50712 35692 50764 35698
rect 50712 35634 50764 35640
rect 50160 35488 50212 35494
rect 50160 35430 50212 35436
rect 50620 35488 50672 35494
rect 50620 35430 50672 35436
rect 50172 35086 50200 35430
rect 49976 35080 50028 35086
rect 49882 35048 49938 35057
rect 49976 35022 50028 35028
rect 50160 35080 50212 35086
rect 50160 35022 50212 35028
rect 49882 34983 49938 34992
rect 49896 34746 49924 34983
rect 49988 34746 50016 35022
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 49884 34740 49936 34746
rect 49884 34682 49936 34688
rect 49976 34740 50028 34746
rect 49976 34682 50028 34688
rect 50252 34672 50304 34678
rect 50250 34640 50252 34649
rect 50304 34640 50306 34649
rect 49884 34604 49936 34610
rect 50160 34604 50212 34610
rect 49884 34546 49936 34552
rect 49988 34564 50160 34592
rect 49896 33998 49924 34546
rect 49884 33992 49936 33998
rect 49988 33969 50016 34564
rect 50250 34575 50306 34584
rect 50160 34546 50212 34552
rect 50068 33992 50120 33998
rect 49884 33934 49936 33940
rect 49974 33960 50030 33969
rect 50068 33934 50120 33940
rect 49974 33895 50030 33904
rect 49988 33590 50016 33895
rect 49976 33584 50028 33590
rect 49976 33526 50028 33532
rect 50080 32978 50108 33934
rect 50160 33924 50212 33930
rect 50160 33866 50212 33872
rect 50172 33114 50200 33866
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50632 33658 50660 35430
rect 50724 34626 50752 35634
rect 50804 34672 50856 34678
rect 50724 34620 50804 34626
rect 50724 34614 50856 34620
rect 50724 34598 50844 34614
rect 50804 34400 50856 34406
rect 50804 34342 50856 34348
rect 50620 33652 50672 33658
rect 50620 33594 50672 33600
rect 50816 33454 50844 34342
rect 50908 33998 50936 38950
rect 51080 38412 51132 38418
rect 51080 38354 51132 38360
rect 50988 34740 51040 34746
rect 50988 34682 51040 34688
rect 50896 33992 50948 33998
rect 50896 33934 50948 33940
rect 50908 33590 50936 33934
rect 50896 33584 50948 33590
rect 50896 33526 50948 33532
rect 51000 33454 51028 34682
rect 51092 34490 51120 38354
rect 51184 35766 51212 39238
rect 51276 37330 51304 40326
rect 51356 39976 51408 39982
rect 51356 39918 51408 39924
rect 51264 37324 51316 37330
rect 51264 37266 51316 37272
rect 51172 35760 51224 35766
rect 51172 35702 51224 35708
rect 51184 35222 51212 35702
rect 51172 35216 51224 35222
rect 51172 35158 51224 35164
rect 51264 35148 51316 35154
rect 51264 35090 51316 35096
rect 51172 34944 51224 34950
rect 51172 34886 51224 34892
rect 51184 34610 51212 34886
rect 51172 34604 51224 34610
rect 51172 34546 51224 34552
rect 51092 34462 51212 34490
rect 51080 34400 51132 34406
rect 51080 34342 51132 34348
rect 51092 33522 51120 34342
rect 51080 33516 51132 33522
rect 51080 33458 51132 33464
rect 50804 33448 50856 33454
rect 50804 33390 50856 33396
rect 50988 33448 51040 33454
rect 50988 33390 51040 33396
rect 51080 33380 51132 33386
rect 51080 33322 51132 33328
rect 50160 33108 50212 33114
rect 50160 33050 50212 33056
rect 50068 32972 50120 32978
rect 50068 32914 50120 32920
rect 50172 32842 50200 33050
rect 51092 32842 51120 33322
rect 50160 32836 50212 32842
rect 50160 32778 50212 32784
rect 50896 32836 50948 32842
rect 50896 32778 50948 32784
rect 51080 32836 51132 32842
rect 51080 32778 51132 32784
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 50908 32434 50936 32778
rect 50068 32428 50120 32434
rect 50068 32370 50120 32376
rect 50896 32428 50948 32434
rect 50896 32370 50948 32376
rect 49974 32328 50030 32337
rect 49974 32263 49976 32272
rect 50028 32263 50030 32272
rect 49976 32234 50028 32240
rect 50080 31754 50108 32370
rect 50908 31822 50936 32370
rect 50896 31816 50948 31822
rect 50896 31758 50948 31764
rect 51080 31816 51132 31822
rect 51080 31758 51132 31764
rect 49804 31726 49924 31754
rect 49700 31476 49752 31482
rect 49700 31418 49752 31424
rect 49332 31340 49384 31346
rect 49332 31282 49384 31288
rect 49516 31340 49568 31346
rect 49516 31282 49568 31288
rect 49240 31272 49292 31278
rect 49240 31214 49292 31220
rect 49148 30932 49200 30938
rect 49148 30874 49200 30880
rect 48780 30864 48832 30870
rect 48780 30806 48832 30812
rect 48872 30728 48924 30734
rect 48872 30670 48924 30676
rect 48688 30252 48740 30258
rect 48688 30194 48740 30200
rect 48700 29238 48728 30194
rect 48780 29708 48832 29714
rect 48780 29650 48832 29656
rect 48688 29232 48740 29238
rect 48688 29174 48740 29180
rect 48504 28960 48556 28966
rect 48504 28902 48556 28908
rect 48792 28762 48820 29650
rect 47952 28756 48004 28762
rect 47952 28698 48004 28704
rect 48780 28756 48832 28762
rect 48780 28698 48832 28704
rect 47964 28626 47992 28698
rect 47952 28620 48004 28626
rect 47952 28562 48004 28568
rect 47768 28552 47820 28558
rect 47768 28494 47820 28500
rect 47860 28552 47912 28558
rect 47860 28494 47912 28500
rect 47780 27878 47808 28494
rect 47872 28150 47900 28494
rect 47964 28218 47992 28562
rect 48042 28384 48098 28393
rect 48042 28319 48098 28328
rect 47952 28212 48004 28218
rect 47952 28154 48004 28160
rect 47860 28144 47912 28150
rect 47860 28086 47912 28092
rect 47768 27872 47820 27878
rect 47768 27814 47820 27820
rect 47780 27674 47808 27814
rect 47872 27674 47900 28086
rect 48056 28082 48084 28319
rect 48320 28212 48372 28218
rect 48320 28154 48372 28160
rect 48044 28076 48096 28082
rect 48044 28018 48096 28024
rect 47768 27668 47820 27674
rect 47768 27610 47820 27616
rect 47860 27668 47912 27674
rect 47860 27610 47912 27616
rect 47676 27532 47728 27538
rect 47676 27474 47728 27480
rect 47308 27464 47360 27470
rect 47308 27406 47360 27412
rect 47320 27062 47348 27406
rect 47308 27056 47360 27062
rect 47308 26998 47360 27004
rect 47688 26790 47716 27474
rect 48332 27470 48360 28154
rect 48884 28082 48912 30670
rect 49160 30394 49188 30874
rect 49148 30388 49200 30394
rect 49148 30330 49200 30336
rect 49252 30258 49280 31214
rect 49344 30326 49372 31282
rect 49332 30320 49384 30326
rect 49332 30262 49384 30268
rect 49528 30258 49556 31282
rect 49712 30734 49740 31418
rect 49700 30728 49752 30734
rect 49700 30670 49752 30676
rect 49240 30252 49292 30258
rect 49240 30194 49292 30200
rect 49516 30252 49568 30258
rect 49516 30194 49568 30200
rect 49528 30122 49556 30194
rect 49516 30116 49568 30122
rect 49516 30058 49568 30064
rect 49608 30116 49660 30122
rect 49608 30058 49660 30064
rect 49424 29232 49476 29238
rect 49424 29174 49476 29180
rect 48872 28076 48924 28082
rect 48872 28018 48924 28024
rect 48964 27940 49016 27946
rect 48964 27882 49016 27888
rect 48872 27600 48924 27606
rect 48872 27542 48924 27548
rect 48136 27464 48188 27470
rect 48136 27406 48188 27412
rect 48320 27464 48372 27470
rect 48320 27406 48372 27412
rect 48148 27130 48176 27406
rect 48136 27124 48188 27130
rect 48136 27066 48188 27072
rect 48044 26988 48096 26994
rect 48044 26930 48096 26936
rect 47676 26784 47728 26790
rect 47676 26726 47728 26732
rect 47124 26580 47176 26586
rect 47124 26522 47176 26528
rect 47216 26580 47268 26586
rect 47216 26522 47268 26528
rect 48056 26246 48084 26930
rect 47676 26240 47728 26246
rect 47676 26182 47728 26188
rect 48044 26240 48096 26246
rect 48044 26182 48096 26188
rect 47688 25362 47716 26182
rect 48884 25906 48912 27542
rect 48976 27062 49004 27882
rect 49436 27470 49464 29174
rect 49620 28218 49648 30058
rect 49896 29510 49924 31726
rect 49976 31748 50108 31754
rect 50028 31726 50108 31748
rect 49976 31690 50028 31696
rect 49988 31278 50016 31690
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50712 31408 50764 31414
rect 50712 31350 50764 31356
rect 49976 31272 50028 31278
rect 49976 31214 50028 31220
rect 49988 30190 50016 31214
rect 50724 30938 50752 31350
rect 50908 31346 50936 31758
rect 51092 31346 51120 31758
rect 51184 31414 51212 34462
rect 51276 33046 51304 35090
rect 51368 34202 51396 39918
rect 51448 38752 51500 38758
rect 51448 38694 51500 38700
rect 51460 38282 51488 38694
rect 51552 38282 51580 40598
rect 51644 40594 51672 40870
rect 51632 40588 51684 40594
rect 51632 40530 51684 40536
rect 51908 40384 51960 40390
rect 51908 40326 51960 40332
rect 51920 40050 51948 40326
rect 51724 40044 51776 40050
rect 51724 39986 51776 39992
rect 51908 40044 51960 40050
rect 51908 39986 51960 39992
rect 51632 39432 51684 39438
rect 51632 39374 51684 39380
rect 51644 38554 51672 39374
rect 51736 38758 51764 39986
rect 52104 39098 52132 44202
rect 52656 43994 52684 44270
rect 53104 44192 53156 44198
rect 53104 44134 53156 44140
rect 52644 43988 52696 43994
rect 52644 43930 52696 43936
rect 52276 43784 52328 43790
rect 52276 43726 52328 43732
rect 52920 43784 52972 43790
rect 52920 43726 52972 43732
rect 52288 43314 52316 43726
rect 52932 43314 52960 43726
rect 53116 43314 53144 44134
rect 53852 43994 53880 44270
rect 54484 44192 54536 44198
rect 54484 44134 54536 44140
rect 53840 43988 53892 43994
rect 53840 43930 53892 43936
rect 54496 43790 54524 44134
rect 55140 43994 55168 44406
rect 55404 44396 55456 44402
rect 55404 44338 55456 44344
rect 55312 44328 55364 44334
rect 55312 44270 55364 44276
rect 55128 43988 55180 43994
rect 55128 43930 55180 43936
rect 53840 43784 53892 43790
rect 53840 43726 53892 43732
rect 54300 43784 54352 43790
rect 54300 43726 54352 43732
rect 54484 43784 54536 43790
rect 54484 43726 54536 43732
rect 52276 43308 52328 43314
rect 52276 43250 52328 43256
rect 52920 43308 52972 43314
rect 52920 43250 52972 43256
rect 53104 43308 53156 43314
rect 53104 43250 53156 43256
rect 53472 43308 53524 43314
rect 53472 43250 53524 43256
rect 52288 42362 52316 43250
rect 52932 42906 52960 43250
rect 52920 42900 52972 42906
rect 52920 42842 52972 42848
rect 53116 42634 53144 43250
rect 53484 42702 53512 43250
rect 53852 42770 53880 43726
rect 54312 43450 54340 43726
rect 54760 43648 54812 43654
rect 54760 43590 54812 43596
rect 54300 43444 54352 43450
rect 54300 43386 54352 43392
rect 54024 43308 54076 43314
rect 54024 43250 54076 43256
rect 54392 43308 54444 43314
rect 54392 43250 54444 43256
rect 53840 42764 53892 42770
rect 53840 42706 53892 42712
rect 53472 42696 53524 42702
rect 53472 42638 53524 42644
rect 53104 42628 53156 42634
rect 53104 42570 53156 42576
rect 52276 42356 52328 42362
rect 52276 42298 52328 42304
rect 52552 41540 52604 41546
rect 52552 41482 52604 41488
rect 52184 41132 52236 41138
rect 52184 41074 52236 41080
rect 52196 40458 52224 41074
rect 52460 41064 52512 41070
rect 52460 41006 52512 41012
rect 52472 40730 52500 41006
rect 52460 40724 52512 40730
rect 52460 40666 52512 40672
rect 52184 40452 52236 40458
rect 52184 40394 52236 40400
rect 52472 40390 52500 40666
rect 52460 40384 52512 40390
rect 52460 40326 52512 40332
rect 52092 39092 52144 39098
rect 52092 39034 52144 39040
rect 52184 38956 52236 38962
rect 52184 38898 52236 38904
rect 51908 38888 51960 38894
rect 51908 38830 51960 38836
rect 51724 38752 51776 38758
rect 51724 38694 51776 38700
rect 51632 38548 51684 38554
rect 51632 38490 51684 38496
rect 51448 38276 51500 38282
rect 51448 38218 51500 38224
rect 51540 38276 51592 38282
rect 51540 38218 51592 38224
rect 51460 35816 51488 38218
rect 51460 35788 51580 35816
rect 51448 35692 51500 35698
rect 51448 35634 51500 35640
rect 51460 34649 51488 35634
rect 51446 34640 51502 34649
rect 51446 34575 51448 34584
rect 51500 34575 51502 34584
rect 51448 34546 51500 34552
rect 51460 34515 51488 34546
rect 51356 34196 51408 34202
rect 51356 34138 51408 34144
rect 51368 33862 51396 34138
rect 51356 33856 51408 33862
rect 51356 33798 51408 33804
rect 51356 33516 51408 33522
rect 51356 33458 51408 33464
rect 51368 33114 51396 33458
rect 51356 33108 51408 33114
rect 51356 33050 51408 33056
rect 51264 33040 51316 33046
rect 51264 32982 51316 32988
rect 51276 32434 51304 32982
rect 51552 32502 51580 35788
rect 51644 35630 51672 38490
rect 51920 37942 51948 38830
rect 52196 38554 52224 38898
rect 52184 38548 52236 38554
rect 52184 38490 52236 38496
rect 52196 38010 52224 38490
rect 52184 38004 52236 38010
rect 52184 37946 52236 37952
rect 51908 37936 51960 37942
rect 51908 37878 51960 37884
rect 51816 37324 51868 37330
rect 51816 37266 51868 37272
rect 51632 35624 51684 35630
rect 51632 35566 51684 35572
rect 51644 34202 51672 35566
rect 51722 35048 51778 35057
rect 51722 34983 51778 34992
rect 51736 34746 51764 34983
rect 51724 34740 51776 34746
rect 51724 34682 51776 34688
rect 51724 34604 51776 34610
rect 51724 34546 51776 34552
rect 51632 34196 51684 34202
rect 51632 34138 51684 34144
rect 51644 34066 51672 34138
rect 51632 34060 51684 34066
rect 51632 34002 51684 34008
rect 51736 33862 51764 34546
rect 51724 33856 51776 33862
rect 51724 33798 51776 33804
rect 51828 33674 51856 37266
rect 51736 33646 51856 33674
rect 51540 32496 51592 32502
rect 51540 32438 51592 32444
rect 51264 32428 51316 32434
rect 51264 32370 51316 32376
rect 51356 31680 51408 31686
rect 51356 31622 51408 31628
rect 51264 31476 51316 31482
rect 51264 31418 51316 31424
rect 51172 31408 51224 31414
rect 51172 31350 51224 31356
rect 50896 31340 50948 31346
rect 50896 31282 50948 31288
rect 51080 31340 51132 31346
rect 51080 31282 51132 31288
rect 50712 30932 50764 30938
rect 50712 30874 50764 30880
rect 51092 30802 51120 31282
rect 51184 31142 51212 31350
rect 51172 31136 51224 31142
rect 51172 31078 51224 31084
rect 51080 30796 51132 30802
rect 51080 30738 51132 30744
rect 51172 30728 51224 30734
rect 51172 30670 51224 30676
rect 50988 30660 51040 30666
rect 50988 30602 51040 30608
rect 50160 30592 50212 30598
rect 50160 30534 50212 30540
rect 49976 30184 50028 30190
rect 49976 30126 50028 30132
rect 49884 29504 49936 29510
rect 49804 29464 49884 29492
rect 49804 29170 49832 29464
rect 49884 29446 49936 29452
rect 49988 29306 50016 30126
rect 50172 29782 50200 30534
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 51000 30326 51028 30602
rect 50988 30320 51040 30326
rect 50988 30262 51040 30268
rect 50804 30184 50856 30190
rect 50804 30126 50856 30132
rect 50160 29776 50212 29782
rect 50160 29718 50212 29724
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 49976 29300 50028 29306
rect 49976 29242 50028 29248
rect 50620 29300 50672 29306
rect 50620 29242 50672 29248
rect 49792 29164 49844 29170
rect 49792 29106 49844 29112
rect 49884 29164 49936 29170
rect 49884 29106 49936 29112
rect 49608 28212 49660 28218
rect 49608 28154 49660 28160
rect 49896 28082 49924 29106
rect 50068 29096 50120 29102
rect 50068 29038 50120 29044
rect 50080 28218 50108 29038
rect 50632 29034 50660 29242
rect 50620 29028 50672 29034
rect 50620 28970 50672 28976
rect 50632 28558 50660 28970
rect 50160 28552 50212 28558
rect 50160 28494 50212 28500
rect 50620 28552 50672 28558
rect 50620 28494 50672 28500
rect 50068 28212 50120 28218
rect 50068 28154 50120 28160
rect 49884 28076 49936 28082
rect 49884 28018 49936 28024
rect 49608 27940 49660 27946
rect 49608 27882 49660 27888
rect 49424 27464 49476 27470
rect 49424 27406 49476 27412
rect 49620 27402 49648 27882
rect 49896 27538 49924 28018
rect 50068 28008 50120 28014
rect 50068 27950 50120 27956
rect 49884 27532 49936 27538
rect 49884 27474 49936 27480
rect 49240 27396 49292 27402
rect 49240 27338 49292 27344
rect 49608 27396 49660 27402
rect 49608 27338 49660 27344
rect 48964 27056 49016 27062
rect 48964 26998 49016 27004
rect 48976 26382 49004 26998
rect 49252 26858 49280 27338
rect 49332 27124 49384 27130
rect 49332 27066 49384 27072
rect 49240 26852 49292 26858
rect 49240 26794 49292 26800
rect 49344 26790 49372 27066
rect 49896 27062 49924 27474
rect 49884 27056 49936 27062
rect 49884 26998 49936 27004
rect 49700 26920 49752 26926
rect 49700 26862 49752 26868
rect 49332 26784 49384 26790
rect 49332 26726 49384 26732
rect 48964 26376 49016 26382
rect 48964 26318 49016 26324
rect 49240 26036 49292 26042
rect 49240 25978 49292 25984
rect 48872 25900 48924 25906
rect 48872 25842 48924 25848
rect 47768 25696 47820 25702
rect 47768 25638 47820 25644
rect 47676 25356 47728 25362
rect 47676 25298 47728 25304
rect 47780 25294 47808 25638
rect 48884 25294 48912 25842
rect 49252 25702 49280 25978
rect 49712 25906 49740 26862
rect 49896 26314 49924 26998
rect 50080 26840 50108 27950
rect 50172 27334 50200 28494
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50160 27328 50212 27334
rect 50160 27270 50212 27276
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50344 26920 50396 26926
rect 50344 26862 50396 26868
rect 50160 26852 50212 26858
rect 50080 26812 50160 26840
rect 50160 26794 50212 26800
rect 50172 26586 50200 26794
rect 50356 26790 50384 26862
rect 50344 26784 50396 26790
rect 50344 26726 50396 26732
rect 50160 26580 50212 26586
rect 50160 26522 50212 26528
rect 50172 26382 50200 26522
rect 50356 26382 50384 26726
rect 50632 26382 50660 28494
rect 50816 27402 50844 30126
rect 51000 29306 51028 30262
rect 51184 29646 51212 30670
rect 51276 30258 51304 31418
rect 51368 30938 51396 31622
rect 51356 30932 51408 30938
rect 51356 30874 51408 30880
rect 51264 30252 51316 30258
rect 51264 30194 51316 30200
rect 51172 29640 51224 29646
rect 51172 29582 51224 29588
rect 51448 29640 51500 29646
rect 51448 29582 51500 29588
rect 50988 29300 51040 29306
rect 50988 29242 51040 29248
rect 51000 29102 51028 29242
rect 50988 29096 51040 29102
rect 50988 29038 51040 29044
rect 51080 28076 51132 28082
rect 51080 28018 51132 28024
rect 50804 27396 50856 27402
rect 50804 27338 50856 27344
rect 50712 26920 50764 26926
rect 50712 26862 50764 26868
rect 50724 26518 50752 26862
rect 51092 26858 51120 28018
rect 51184 27402 51212 29582
rect 51460 29170 51488 29582
rect 51736 29288 51764 33646
rect 51816 33040 51868 33046
rect 51816 32982 51868 32988
rect 51828 32502 51856 32982
rect 51816 32496 51868 32502
rect 51816 32438 51868 32444
rect 51920 31210 51948 37878
rect 52184 37868 52236 37874
rect 52184 37810 52236 37816
rect 52196 37126 52224 37810
rect 52184 37120 52236 37126
rect 52184 37062 52236 37068
rect 52276 36576 52328 36582
rect 52276 36518 52328 36524
rect 52288 36242 52316 36518
rect 52276 36236 52328 36242
rect 52276 36178 52328 36184
rect 52368 36168 52420 36174
rect 52368 36110 52420 36116
rect 52092 36100 52144 36106
rect 52092 36042 52144 36048
rect 52104 35290 52132 36042
rect 52380 35290 52408 36110
rect 52092 35284 52144 35290
rect 52092 35226 52144 35232
rect 52368 35284 52420 35290
rect 52368 35226 52420 35232
rect 52276 35216 52328 35222
rect 52276 35158 52328 35164
rect 52288 34746 52316 35158
rect 52472 35086 52500 40326
rect 52564 35154 52592 41482
rect 52736 40996 52788 41002
rect 52736 40938 52788 40944
rect 52748 40526 52776 40938
rect 52736 40520 52788 40526
rect 52736 40462 52788 40468
rect 52748 40186 52776 40462
rect 52736 40180 52788 40186
rect 52736 40122 52788 40128
rect 52828 40180 52880 40186
rect 52828 40122 52880 40128
rect 52552 35148 52604 35154
rect 52552 35090 52604 35096
rect 52460 35080 52512 35086
rect 52460 35022 52512 35028
rect 52460 34944 52512 34950
rect 52460 34886 52512 34892
rect 52276 34740 52328 34746
rect 52276 34682 52328 34688
rect 52000 34604 52052 34610
rect 52000 34546 52052 34552
rect 52184 34604 52236 34610
rect 52184 34546 52236 34552
rect 52012 33658 52040 34546
rect 52196 33930 52224 34546
rect 52472 33998 52500 34886
rect 52564 34066 52592 35090
rect 52644 35080 52696 35086
rect 52644 35022 52696 35028
rect 52656 34202 52684 35022
rect 52748 34950 52776 40122
rect 52840 39914 52868 40122
rect 52828 39908 52880 39914
rect 52828 39850 52880 39856
rect 53196 39840 53248 39846
rect 53196 39782 53248 39788
rect 53012 38344 53064 38350
rect 53012 38286 53064 38292
rect 52736 34944 52788 34950
rect 52736 34886 52788 34892
rect 52644 34196 52696 34202
rect 52644 34138 52696 34144
rect 52552 34060 52604 34066
rect 52552 34002 52604 34008
rect 52736 34060 52788 34066
rect 52736 34002 52788 34008
rect 52368 33992 52420 33998
rect 52368 33934 52420 33940
rect 52460 33992 52512 33998
rect 52460 33934 52512 33940
rect 52184 33924 52236 33930
rect 52184 33866 52236 33872
rect 52000 33652 52052 33658
rect 52000 33594 52052 33600
rect 52196 31754 52224 33866
rect 52380 33590 52408 33934
rect 52368 33584 52420 33590
rect 52368 33526 52420 33532
rect 52644 32428 52696 32434
rect 52644 32370 52696 32376
rect 52552 32360 52604 32366
rect 52552 32302 52604 32308
rect 52564 31822 52592 32302
rect 52656 31822 52684 32370
rect 52552 31816 52604 31822
rect 52552 31758 52604 31764
rect 52644 31816 52696 31822
rect 52644 31758 52696 31764
rect 52104 31726 52224 31754
rect 52104 31362 52132 31726
rect 52184 31408 52236 31414
rect 52104 31356 52184 31362
rect 52104 31350 52236 31356
rect 52000 31340 52052 31346
rect 52000 31282 52052 31288
rect 52104 31334 52224 31350
rect 52368 31340 52420 31346
rect 51908 31204 51960 31210
rect 51908 31146 51960 31152
rect 52012 30122 52040 31282
rect 52104 30666 52132 31334
rect 52368 31282 52420 31288
rect 52380 30666 52408 31282
rect 52656 30938 52684 31758
rect 52644 30932 52696 30938
rect 52644 30874 52696 30880
rect 52092 30660 52144 30666
rect 52368 30660 52420 30666
rect 52092 30602 52144 30608
rect 52288 30620 52368 30648
rect 52104 30258 52132 30602
rect 52092 30252 52144 30258
rect 52092 30194 52144 30200
rect 52000 30116 52052 30122
rect 52000 30058 52052 30064
rect 51816 29300 51868 29306
rect 51736 29260 51816 29288
rect 51816 29242 51868 29248
rect 51448 29164 51500 29170
rect 51448 29106 51500 29112
rect 51908 28552 51960 28558
rect 51908 28494 51960 28500
rect 51632 28484 51684 28490
rect 51632 28426 51684 28432
rect 51644 28082 51672 28426
rect 51632 28076 51684 28082
rect 51632 28018 51684 28024
rect 51356 28008 51408 28014
rect 51356 27950 51408 27956
rect 51172 27396 51224 27402
rect 51172 27338 51224 27344
rect 51368 27130 51396 27950
rect 51448 27464 51500 27470
rect 51448 27406 51500 27412
rect 51356 27124 51408 27130
rect 51356 27066 51408 27072
rect 51460 26926 51488 27406
rect 51540 27328 51592 27334
rect 51540 27270 51592 27276
rect 51552 27130 51580 27270
rect 51540 27124 51592 27130
rect 51540 27066 51592 27072
rect 51644 27062 51672 28018
rect 51920 27946 51948 28494
rect 51908 27940 51960 27946
rect 51908 27882 51960 27888
rect 51920 27130 51948 27882
rect 51908 27124 51960 27130
rect 51908 27066 51960 27072
rect 51632 27056 51684 27062
rect 51632 26998 51684 27004
rect 51448 26920 51500 26926
rect 51448 26862 51500 26868
rect 51080 26852 51132 26858
rect 51080 26794 51132 26800
rect 50712 26512 50764 26518
rect 50712 26454 50764 26460
rect 51092 26450 51120 26794
rect 51644 26586 51672 26998
rect 51632 26580 51684 26586
rect 51632 26522 51684 26528
rect 51080 26444 51132 26450
rect 51080 26386 51132 26392
rect 50160 26376 50212 26382
rect 50160 26318 50212 26324
rect 50344 26376 50396 26382
rect 50344 26318 50396 26324
rect 50620 26376 50672 26382
rect 50620 26318 50672 26324
rect 52288 26314 52316 30620
rect 52368 30602 52420 30608
rect 52748 29850 52776 34002
rect 52828 32292 52880 32298
rect 52828 32234 52880 32240
rect 52840 31890 52868 32234
rect 52828 31884 52880 31890
rect 52828 31826 52880 31832
rect 52840 31210 52868 31826
rect 53024 31482 53052 38286
rect 53208 37806 53236 39782
rect 53484 39098 53512 42638
rect 54036 42634 54064 43250
rect 54116 43172 54168 43178
rect 54116 43114 54168 43120
rect 54024 42628 54076 42634
rect 54024 42570 54076 42576
rect 54036 42362 54064 42570
rect 54024 42356 54076 42362
rect 54024 42298 54076 42304
rect 54128 42226 54156 43114
rect 54404 42634 54432 43250
rect 54772 42838 54800 43590
rect 55140 43450 55168 43930
rect 55324 43722 55352 44270
rect 55312 43716 55364 43722
rect 55312 43658 55364 43664
rect 55416 43654 55444 44338
rect 55404 43648 55456 43654
rect 55404 43590 55456 43596
rect 55128 43444 55180 43450
rect 55128 43386 55180 43392
rect 55312 43308 55364 43314
rect 55312 43250 55364 43256
rect 54760 42832 54812 42838
rect 54760 42774 54812 42780
rect 55324 42634 55352 43250
rect 55416 42906 55444 43590
rect 55588 43444 55640 43450
rect 55588 43386 55640 43392
rect 55496 43308 55548 43314
rect 55496 43250 55548 43256
rect 55404 42900 55456 42906
rect 55404 42842 55456 42848
rect 55508 42634 55536 43250
rect 55600 42702 55628 43386
rect 55588 42696 55640 42702
rect 55588 42638 55640 42644
rect 54392 42628 54444 42634
rect 54392 42570 54444 42576
rect 55312 42628 55364 42634
rect 55312 42570 55364 42576
rect 55496 42628 55548 42634
rect 55496 42570 55548 42576
rect 54116 42220 54168 42226
rect 54116 42162 54168 42168
rect 55128 42220 55180 42226
rect 55128 42162 55180 42168
rect 54128 42022 54156 42162
rect 54116 42016 54168 42022
rect 54116 41958 54168 41964
rect 54760 40452 54812 40458
rect 54760 40394 54812 40400
rect 54772 40050 54800 40394
rect 54116 40044 54168 40050
rect 54116 39986 54168 39992
rect 54760 40044 54812 40050
rect 54760 39986 54812 39992
rect 53930 39944 53986 39953
rect 53930 39879 53932 39888
rect 53984 39879 53986 39888
rect 53932 39850 53984 39856
rect 54128 39642 54156 39986
rect 55140 39982 55168 42162
rect 55324 41274 55352 42570
rect 55600 42362 55628 42638
rect 55588 42356 55640 42362
rect 55588 42298 55640 42304
rect 55312 41268 55364 41274
rect 55312 41210 55364 41216
rect 55496 40520 55548 40526
rect 55496 40462 55548 40468
rect 55312 40384 55364 40390
rect 55312 40326 55364 40332
rect 55324 40050 55352 40326
rect 55220 40044 55272 40050
rect 55220 39986 55272 39992
rect 55312 40044 55364 40050
rect 55312 39986 55364 39992
rect 55128 39976 55180 39982
rect 55128 39918 55180 39924
rect 54116 39636 54168 39642
rect 54116 39578 54168 39584
rect 55232 39574 55260 39986
rect 55508 39642 55536 40462
rect 55496 39636 55548 39642
rect 55496 39578 55548 39584
rect 55220 39568 55272 39574
rect 55220 39510 55272 39516
rect 54484 39500 54536 39506
rect 54484 39442 54536 39448
rect 53656 39432 53708 39438
rect 53656 39374 53708 39380
rect 53472 39092 53524 39098
rect 53472 39034 53524 39040
rect 53288 38956 53340 38962
rect 53288 38898 53340 38904
rect 53300 38554 53328 38898
rect 53668 38894 53696 39374
rect 53656 38888 53708 38894
rect 53656 38830 53708 38836
rect 53668 38554 53696 38830
rect 53288 38548 53340 38554
rect 53288 38490 53340 38496
rect 53656 38548 53708 38554
rect 53656 38490 53708 38496
rect 53748 38412 53800 38418
rect 53748 38354 53800 38360
rect 53196 37800 53248 37806
rect 53196 37742 53248 37748
rect 53380 35488 53432 35494
rect 53380 35430 53432 35436
rect 53392 35086 53420 35430
rect 53380 35080 53432 35086
rect 53380 35022 53432 35028
rect 53472 34944 53524 34950
rect 53472 34886 53524 34892
rect 53484 34066 53512 34886
rect 53656 34536 53708 34542
rect 53656 34478 53708 34484
rect 53472 34060 53524 34066
rect 53472 34002 53524 34008
rect 53564 32428 53616 32434
rect 53564 32370 53616 32376
rect 53104 32360 53156 32366
rect 53104 32302 53156 32308
rect 53116 32026 53144 32302
rect 53576 32026 53604 32370
rect 53104 32020 53156 32026
rect 53104 31962 53156 31968
rect 53564 32020 53616 32026
rect 53564 31962 53616 31968
rect 53472 31816 53524 31822
rect 53472 31758 53524 31764
rect 53012 31476 53064 31482
rect 53012 31418 53064 31424
rect 53484 31346 53512 31758
rect 53576 31346 53604 31962
rect 53472 31340 53524 31346
rect 53472 31282 53524 31288
rect 53564 31340 53616 31346
rect 53564 31282 53616 31288
rect 52828 31204 52880 31210
rect 52828 31146 52880 31152
rect 52736 29844 52788 29850
rect 52736 29786 52788 29792
rect 52460 29572 52512 29578
rect 52460 29514 52512 29520
rect 52472 29238 52500 29514
rect 53012 29504 53064 29510
rect 53012 29446 53064 29452
rect 52460 29232 52512 29238
rect 52460 29174 52512 29180
rect 52472 28558 52500 29174
rect 53024 29102 53052 29446
rect 52920 29096 52972 29102
rect 52920 29038 52972 29044
rect 53012 29096 53064 29102
rect 53012 29038 53064 29044
rect 52828 29028 52880 29034
rect 52828 28970 52880 28976
rect 52840 28762 52868 28970
rect 52828 28756 52880 28762
rect 52828 28698 52880 28704
rect 52460 28552 52512 28558
rect 52460 28494 52512 28500
rect 52368 28416 52420 28422
rect 52368 28358 52420 28364
rect 52380 28014 52408 28358
rect 52368 28008 52420 28014
rect 52368 27950 52420 27956
rect 52380 27470 52408 27950
rect 52472 27878 52500 28494
rect 52840 28082 52868 28698
rect 52932 28642 52960 29038
rect 53024 28762 53052 29038
rect 53012 28756 53064 28762
rect 53012 28698 53064 28704
rect 52932 28614 53052 28642
rect 52920 28552 52972 28558
rect 52920 28494 52972 28500
rect 52828 28076 52880 28082
rect 52828 28018 52880 28024
rect 52460 27872 52512 27878
rect 52460 27814 52512 27820
rect 52368 27464 52420 27470
rect 52368 27406 52420 27412
rect 52472 26790 52500 27814
rect 52932 27674 52960 28494
rect 53024 28218 53052 28614
rect 53196 28484 53248 28490
rect 53196 28426 53248 28432
rect 53012 28212 53064 28218
rect 53012 28154 53064 28160
rect 52920 27668 52972 27674
rect 52920 27610 52972 27616
rect 53024 27538 53052 28154
rect 53104 28008 53156 28014
rect 53104 27950 53156 27956
rect 53116 27878 53144 27950
rect 53104 27872 53156 27878
rect 53104 27814 53156 27820
rect 53012 27532 53064 27538
rect 53012 27474 53064 27480
rect 53208 27470 53236 28426
rect 53484 28218 53512 31282
rect 53668 31210 53696 34478
rect 53760 32570 53788 38354
rect 53932 37732 53984 37738
rect 53932 37674 53984 37680
rect 53944 36718 53972 37674
rect 54024 36780 54076 36786
rect 54024 36722 54076 36728
rect 53932 36712 53984 36718
rect 53932 36654 53984 36660
rect 53932 33584 53984 33590
rect 53932 33526 53984 33532
rect 53944 32774 53972 33526
rect 53932 32768 53984 32774
rect 53932 32710 53984 32716
rect 53748 32564 53800 32570
rect 53748 32506 53800 32512
rect 53748 31816 53800 31822
rect 53748 31758 53800 31764
rect 53760 31414 53788 31758
rect 53748 31408 53800 31414
rect 53748 31350 53800 31356
rect 53656 31204 53708 31210
rect 53656 31146 53708 31152
rect 54036 29850 54064 36722
rect 54496 34202 54524 39442
rect 54944 36712 54996 36718
rect 54944 36654 54996 36660
rect 54956 36378 54984 36654
rect 54944 36372 54996 36378
rect 54944 36314 54996 36320
rect 55588 35012 55640 35018
rect 55588 34954 55640 34960
rect 54484 34196 54536 34202
rect 54484 34138 54536 34144
rect 55600 33998 55628 34954
rect 54484 33992 54536 33998
rect 54484 33934 54536 33940
rect 54668 33992 54720 33998
rect 54668 33934 54720 33940
rect 55588 33992 55640 33998
rect 55588 33934 55640 33940
rect 54208 33584 54260 33590
rect 54208 33526 54260 33532
rect 54116 33312 54168 33318
rect 54116 33254 54168 33260
rect 54128 32910 54156 33254
rect 54116 32904 54168 32910
rect 54116 32846 54168 32852
rect 54220 32842 54248 33526
rect 54496 33114 54524 33934
rect 54680 33386 54708 33934
rect 55496 33856 55548 33862
rect 55496 33798 55548 33804
rect 54760 33516 54812 33522
rect 54760 33458 54812 33464
rect 55404 33516 55456 33522
rect 55404 33458 55456 33464
rect 54668 33380 54720 33386
rect 54668 33322 54720 33328
rect 54484 33108 54536 33114
rect 54484 33050 54536 33056
rect 54772 32910 54800 33458
rect 54576 32904 54628 32910
rect 54576 32846 54628 32852
rect 54760 32904 54812 32910
rect 54760 32846 54812 32852
rect 54208 32836 54260 32842
rect 54208 32778 54260 32784
rect 54588 31482 54616 32846
rect 54668 32292 54720 32298
rect 54668 32234 54720 32240
rect 54576 31476 54628 31482
rect 54576 31418 54628 31424
rect 54680 30734 54708 32234
rect 54772 31958 54800 32846
rect 55416 32026 55444 33458
rect 55508 32842 55536 33798
rect 55600 33658 55628 33934
rect 55588 33652 55640 33658
rect 55588 33594 55640 33600
rect 55588 33108 55640 33114
rect 55588 33050 55640 33056
rect 55496 32836 55548 32842
rect 55496 32778 55548 32784
rect 55508 32434 55536 32778
rect 55496 32428 55548 32434
rect 55496 32370 55548 32376
rect 55600 32366 55628 33050
rect 55588 32360 55640 32366
rect 55588 32302 55640 32308
rect 55404 32020 55456 32026
rect 55404 31962 55456 31968
rect 54760 31952 54812 31958
rect 54760 31894 54812 31900
rect 55600 31482 55628 32302
rect 55404 31476 55456 31482
rect 55404 31418 55456 31424
rect 55588 31476 55640 31482
rect 55588 31418 55640 31424
rect 54668 30728 54720 30734
rect 54668 30670 54720 30676
rect 54208 30592 54260 30598
rect 54208 30534 54260 30540
rect 54220 30326 54248 30534
rect 54208 30320 54260 30326
rect 54208 30262 54260 30268
rect 54024 29844 54076 29850
rect 54024 29786 54076 29792
rect 54024 29708 54076 29714
rect 54024 29650 54076 29656
rect 54036 29102 54064 29650
rect 54220 29646 54248 30262
rect 54680 30258 54708 30670
rect 55416 30666 55444 31418
rect 55588 31204 55640 31210
rect 55588 31146 55640 31152
rect 55600 30734 55628 31146
rect 55588 30728 55640 30734
rect 55588 30670 55640 30676
rect 54760 30660 54812 30666
rect 54760 30602 54812 30608
rect 55404 30660 55456 30666
rect 55404 30602 55456 30608
rect 54772 30258 54800 30602
rect 54668 30252 54720 30258
rect 54668 30194 54720 30200
rect 54760 30252 54812 30258
rect 54760 30194 54812 30200
rect 54208 29640 54260 29646
rect 54208 29582 54260 29588
rect 54392 29504 54444 29510
rect 54392 29446 54444 29452
rect 54404 29306 54432 29446
rect 54772 29306 54800 30194
rect 55416 29850 55444 30602
rect 55404 29844 55456 29850
rect 55404 29786 55456 29792
rect 55312 29640 55364 29646
rect 55312 29582 55364 29588
rect 55496 29640 55548 29646
rect 55496 29582 55548 29588
rect 54392 29300 54444 29306
rect 54392 29242 54444 29248
rect 54760 29300 54812 29306
rect 54760 29242 54812 29248
rect 54024 29096 54076 29102
rect 54024 29038 54076 29044
rect 55324 28762 55352 29582
rect 55312 28756 55364 28762
rect 55312 28698 55364 28704
rect 55220 28688 55272 28694
rect 55220 28630 55272 28636
rect 54668 28552 54720 28558
rect 54668 28494 54720 28500
rect 54392 28484 54444 28490
rect 54392 28426 54444 28432
rect 53472 28212 53524 28218
rect 53472 28154 53524 28160
rect 54404 28064 54432 28426
rect 54680 28082 54708 28494
rect 54484 28076 54536 28082
rect 54404 28036 54484 28064
rect 54484 28018 54536 28024
rect 54668 28076 54720 28082
rect 54668 28018 54720 28024
rect 53656 27872 53708 27878
rect 53656 27814 53708 27820
rect 53668 27470 53696 27814
rect 54496 27538 54524 28018
rect 55232 27985 55260 28630
rect 55508 28218 55536 29582
rect 55496 28212 55548 28218
rect 55496 28154 55548 28160
rect 55218 27976 55274 27985
rect 55218 27911 55274 27920
rect 54484 27532 54536 27538
rect 54484 27474 54536 27480
rect 53196 27464 53248 27470
rect 53196 27406 53248 27412
rect 53656 27464 53708 27470
rect 53656 27406 53708 27412
rect 52460 26784 52512 26790
rect 52460 26726 52512 26732
rect 49884 26308 49936 26314
rect 49884 26250 49936 26256
rect 51264 26308 51316 26314
rect 51264 26250 51316 26256
rect 52276 26308 52328 26314
rect 52276 26250 52328 26256
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 51276 26042 51304 26250
rect 51264 26036 51316 26042
rect 51264 25978 51316 25984
rect 49700 25900 49752 25906
rect 49700 25842 49752 25848
rect 49240 25696 49292 25702
rect 49240 25638 49292 25644
rect 47768 25288 47820 25294
rect 47768 25230 47820 25236
rect 48872 25288 48924 25294
rect 48872 25230 48924 25236
rect 47308 25152 47360 25158
rect 47308 25094 47360 25100
rect 47676 25152 47728 25158
rect 47676 25094 47728 25100
rect 47216 24948 47268 24954
rect 47216 24890 47268 24896
rect 46756 24812 46808 24818
rect 46584 24772 46756 24800
rect 46480 24404 46532 24410
rect 46480 24346 46532 24352
rect 46584 24138 46612 24772
rect 46756 24754 46808 24760
rect 47228 24682 47256 24890
rect 46664 24676 46716 24682
rect 46664 24618 46716 24624
rect 47216 24676 47268 24682
rect 47216 24618 47268 24624
rect 46572 24132 46624 24138
rect 46572 24074 46624 24080
rect 46388 23792 46440 23798
rect 46388 23734 46440 23740
rect 46584 23662 46612 24074
rect 46676 23730 46704 24618
rect 46940 24336 46992 24342
rect 46940 24278 46992 24284
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 46572 23656 46624 23662
rect 46572 23598 46624 23604
rect 46296 23180 46348 23186
rect 46296 23122 46348 23128
rect 46952 23118 46980 24278
rect 47320 24206 47348 25094
rect 47584 24812 47636 24818
rect 47584 24754 47636 24760
rect 47596 24682 47624 24754
rect 47584 24676 47636 24682
rect 47584 24618 47636 24624
rect 47688 24614 47716 25094
rect 47952 24744 48004 24750
rect 47950 24712 47952 24721
rect 48004 24712 48006 24721
rect 49252 24682 49280 25638
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 47950 24647 48006 24656
rect 49240 24676 49292 24682
rect 49240 24618 49292 24624
rect 47676 24608 47728 24614
rect 47676 24550 47728 24556
rect 47952 24268 48004 24274
rect 47952 24210 48004 24216
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 47124 23792 47176 23798
rect 47124 23734 47176 23740
rect 47136 23118 47164 23734
rect 47320 23730 47348 24142
rect 47964 23866 47992 24210
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 47952 23860 48004 23866
rect 47952 23802 48004 23808
rect 47308 23724 47360 23730
rect 47308 23666 47360 23672
rect 47768 23724 47820 23730
rect 47768 23666 47820 23672
rect 47780 23322 47808 23666
rect 47768 23316 47820 23322
rect 47768 23258 47820 23264
rect 46940 23112 46992 23118
rect 46940 23054 46992 23060
rect 47124 23112 47176 23118
rect 47124 23054 47176 23060
rect 45468 22976 45520 22982
rect 45468 22918 45520 22924
rect 45480 22778 45508 22918
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 45468 22772 45520 22778
rect 45468 22714 45520 22720
rect 45192 22636 45244 22642
rect 45192 22578 45244 22584
rect 45204 22234 45232 22578
rect 44640 22228 44692 22234
rect 44640 22170 44692 22176
rect 45192 22228 45244 22234
rect 45192 22170 45244 22176
rect 44272 21888 44324 21894
rect 44272 21830 44324 21836
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 47584 20800 47636 20806
rect 47584 20742 47636 20748
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 46756 19780 46808 19786
rect 46756 19722 46808 19728
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 46768 4078 46796 19722
rect 46756 4072 46808 4078
rect 46756 4014 46808 4020
rect 44548 4004 44600 4010
rect 44548 3946 44600 3952
rect 38476 3936 38528 3942
rect 38476 3878 38528 3884
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 32128 3596 32180 3602
rect 32128 3538 32180 3544
rect 32864 3596 32916 3602
rect 32864 3538 32916 3544
rect 34152 3596 34204 3602
rect 34152 3538 34204 3544
rect 31208 3460 31260 3466
rect 31208 3402 31260 3408
rect 31576 3460 31628 3466
rect 31576 3402 31628 3408
rect 32680 3460 32732 3466
rect 32680 3402 32732 3408
rect 30748 3120 30800 3126
rect 30748 3062 30800 3068
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 30932 2984 30984 2990
rect 30932 2926 30984 2932
rect 28816 2848 28868 2854
rect 28816 2790 28868 2796
rect 30944 800 30972 2926
rect 31116 2848 31168 2854
rect 31116 2790 31168 2796
rect 31128 2446 31156 2790
rect 31220 2650 31248 3402
rect 31208 2644 31260 2650
rect 31208 2586 31260 2592
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31588 800 31616 3402
rect 32692 3194 32720 3402
rect 32680 3188 32732 3194
rect 32680 3130 32732 3136
rect 32876 800 32904 3538
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 38304 3058 38332 3470
rect 38488 3126 38516 3878
rect 43260 3664 43312 3670
rect 43260 3606 43312 3612
rect 43272 3466 43300 3606
rect 43260 3460 43312 3466
rect 43260 3402 43312 3408
rect 44560 3398 44588 3946
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3602 46336 3878
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 44548 3392 44600 3398
rect 44548 3334 44600 3340
rect 38476 3120 38528 3126
rect 38476 3062 38528 3068
rect 46768 3058 46796 4014
rect 47032 3596 47084 3602
rect 47032 3538 47084 3544
rect 46848 3460 46900 3466
rect 46848 3402 46900 3408
rect 46860 3194 46888 3402
rect 46848 3188 46900 3194
rect 46848 3130 46900 3136
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 46756 3052 46808 3058
rect 46756 2994 46808 3000
rect 38660 2984 38712 2990
rect 38660 2926 38712 2932
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 38672 800 38700 2926
rect 47044 800 47072 3538
rect 47596 3058 47624 20742
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 55692 15026 55720 55694
rect 56612 55418 56640 57190
rect 56704 56302 56732 59200
rect 57704 57452 57756 57458
rect 57704 57394 57756 57400
rect 57244 57248 57296 57254
rect 57244 57190 57296 57196
rect 57428 57248 57480 57254
rect 57428 57190 57480 57196
rect 56876 56364 56928 56370
rect 56876 56306 56928 56312
rect 56692 56296 56744 56302
rect 56692 56238 56744 56244
rect 56888 56166 56916 56306
rect 56876 56160 56928 56166
rect 56876 56102 56928 56108
rect 56784 55616 56836 55622
rect 56784 55558 56836 55564
rect 56796 55418 56824 55558
rect 56600 55412 56652 55418
rect 56600 55354 56652 55360
rect 56784 55412 56836 55418
rect 56784 55354 56836 55360
rect 56600 55140 56652 55146
rect 56600 55082 56652 55088
rect 56324 54664 56376 54670
rect 56324 54606 56376 54612
rect 56336 54262 56364 54606
rect 56324 54256 56376 54262
rect 56324 54198 56376 54204
rect 56232 54188 56284 54194
rect 56232 54130 56284 54136
rect 56244 47190 56272 54130
rect 56508 53984 56560 53990
rect 56508 53926 56560 53932
rect 56520 53650 56548 53926
rect 56508 53644 56560 53650
rect 56508 53586 56560 53592
rect 56324 53576 56376 53582
rect 56324 53518 56376 53524
rect 56336 53106 56364 53518
rect 56324 53100 56376 53106
rect 56324 53042 56376 53048
rect 56612 49230 56640 55082
rect 56796 51074 56824 55354
rect 56888 54194 56916 56102
rect 57256 55962 57284 57190
rect 57244 55956 57296 55962
rect 57244 55898 57296 55904
rect 57440 55894 57468 57190
rect 57428 55888 57480 55894
rect 57334 55856 57390 55865
rect 57428 55830 57480 55836
rect 57334 55791 57390 55800
rect 57348 55350 57376 55791
rect 57336 55344 57388 55350
rect 57336 55286 57388 55292
rect 56968 54596 57020 54602
rect 56968 54538 57020 54544
rect 56980 54330 57008 54538
rect 56968 54324 57020 54330
rect 56968 54266 57020 54272
rect 56876 54188 56928 54194
rect 56876 54130 56928 54136
rect 57520 51400 57572 51406
rect 57520 51342 57572 51348
rect 57060 51264 57112 51270
rect 57060 51206 57112 51212
rect 56704 51046 56824 51074
rect 56600 49224 56652 49230
rect 56600 49166 56652 49172
rect 56232 47184 56284 47190
rect 56232 47126 56284 47132
rect 55864 45484 55916 45490
rect 55864 45426 55916 45432
rect 56048 45484 56100 45490
rect 56048 45426 56100 45432
rect 55876 45370 55904 45426
rect 55784 45342 55904 45370
rect 55784 44810 55812 45342
rect 55864 45280 55916 45286
rect 55864 45222 55916 45228
rect 55876 44878 55904 45222
rect 56060 44946 56088 45426
rect 56048 44940 56100 44946
rect 56048 44882 56100 44888
rect 55864 44872 55916 44878
rect 55864 44814 55916 44820
rect 55772 44804 55824 44810
rect 55772 44746 55824 44752
rect 55784 44334 55812 44746
rect 55772 44328 55824 44334
rect 55772 44270 55824 44276
rect 55956 43716 56008 43722
rect 55956 43658 56008 43664
rect 55772 40520 55824 40526
rect 55772 40462 55824 40468
rect 55784 40118 55812 40462
rect 55772 40112 55824 40118
rect 55772 40054 55824 40060
rect 55864 33992 55916 33998
rect 55864 33934 55916 33940
rect 55876 33658 55904 33934
rect 55864 33652 55916 33658
rect 55864 33594 55916 33600
rect 55864 31816 55916 31822
rect 55864 31758 55916 31764
rect 55876 31414 55904 31758
rect 55864 31408 55916 31414
rect 55864 31350 55916 31356
rect 55772 31340 55824 31346
rect 55772 31282 55824 31288
rect 55784 30394 55812 31282
rect 55772 30388 55824 30394
rect 55772 30330 55824 30336
rect 55968 27130 55996 43658
rect 56060 37398 56088 44882
rect 56324 44464 56376 44470
rect 56324 44406 56376 44412
rect 56336 43314 56364 44406
rect 56508 44396 56560 44402
rect 56508 44338 56560 44344
rect 56324 43308 56376 43314
rect 56324 43250 56376 43256
rect 56520 42294 56548 44338
rect 56600 44192 56652 44198
rect 56600 44134 56652 44140
rect 56612 43858 56640 44134
rect 56600 43852 56652 43858
rect 56600 43794 56652 43800
rect 56508 42288 56560 42294
rect 56508 42230 56560 42236
rect 56520 41818 56548 42230
rect 56508 41812 56560 41818
rect 56508 41754 56560 41760
rect 56232 41132 56284 41138
rect 56232 41074 56284 41080
rect 56244 40730 56272 41074
rect 56232 40724 56284 40730
rect 56232 40666 56284 40672
rect 56416 40520 56468 40526
rect 56416 40462 56468 40468
rect 56232 40452 56284 40458
rect 56232 40394 56284 40400
rect 56244 40186 56272 40394
rect 56428 40186 56456 40462
rect 56232 40180 56284 40186
rect 56232 40122 56284 40128
rect 56416 40180 56468 40186
rect 56416 40122 56468 40128
rect 56324 40044 56376 40050
rect 56324 39986 56376 39992
rect 56336 39438 56364 39986
rect 56416 39976 56468 39982
rect 56416 39918 56468 39924
rect 56428 39642 56456 39918
rect 56416 39636 56468 39642
rect 56416 39578 56468 39584
rect 56324 39432 56376 39438
rect 56324 39374 56376 39380
rect 56048 37392 56100 37398
rect 56048 37334 56100 37340
rect 56428 36378 56456 39578
rect 56600 38752 56652 38758
rect 56600 38694 56652 38700
rect 56612 38418 56640 38694
rect 56600 38412 56652 38418
rect 56600 38354 56652 38360
rect 56600 37324 56652 37330
rect 56600 37266 56652 37272
rect 56612 36922 56640 37266
rect 56600 36916 56652 36922
rect 56600 36858 56652 36864
rect 56508 36780 56560 36786
rect 56508 36722 56560 36728
rect 56416 36372 56468 36378
rect 56416 36314 56468 36320
rect 56140 36236 56192 36242
rect 56140 36178 56192 36184
rect 56048 36168 56100 36174
rect 56048 36110 56100 36116
rect 56060 35494 56088 36110
rect 56152 35698 56180 36178
rect 56140 35692 56192 35698
rect 56140 35634 56192 35640
rect 56048 35488 56100 35494
rect 56048 35430 56100 35436
rect 56152 34202 56180 35634
rect 56324 35488 56376 35494
rect 56324 35430 56376 35436
rect 56336 35086 56364 35430
rect 56324 35080 56376 35086
rect 56324 35022 56376 35028
rect 56140 34196 56192 34202
rect 56140 34138 56192 34144
rect 56324 33856 56376 33862
rect 56324 33798 56376 33804
rect 56336 33590 56364 33798
rect 56324 33584 56376 33590
rect 56324 33526 56376 33532
rect 56416 33516 56468 33522
rect 56416 33458 56468 33464
rect 56428 33114 56456 33458
rect 56416 33108 56468 33114
rect 56416 33050 56468 33056
rect 56520 32570 56548 36722
rect 56704 34610 56732 51046
rect 57072 50386 57100 51206
rect 57060 50380 57112 50386
rect 57060 50322 57112 50328
rect 57244 49224 57296 49230
rect 57244 49166 57296 49172
rect 57152 49088 57204 49094
rect 57152 49030 57204 49036
rect 56876 48748 56928 48754
rect 56876 48690 56928 48696
rect 56888 45966 56916 48690
rect 57164 48210 57192 49030
rect 57256 48278 57284 49166
rect 57244 48272 57296 48278
rect 57244 48214 57296 48220
rect 57152 48204 57204 48210
rect 57152 48146 57204 48152
rect 56968 46980 57020 46986
rect 56968 46922 57020 46928
rect 56980 46714 57008 46922
rect 56968 46708 57020 46714
rect 56968 46650 57020 46656
rect 56876 45960 56928 45966
rect 56876 45902 56928 45908
rect 57428 45960 57480 45966
rect 57428 45902 57480 45908
rect 57060 45824 57112 45830
rect 57060 45766 57112 45772
rect 57072 44946 57100 45766
rect 57060 44940 57112 44946
rect 57060 44882 57112 44888
rect 56968 44396 57020 44402
rect 56968 44338 57020 44344
rect 56980 43246 57008 44338
rect 57152 43988 57204 43994
rect 57152 43930 57204 43936
rect 57164 43450 57192 43930
rect 57152 43444 57204 43450
rect 57152 43386 57204 43392
rect 56968 43240 57020 43246
rect 56968 43182 57020 43188
rect 56876 43104 56928 43110
rect 56876 43046 56928 43052
rect 56888 42770 56916 43046
rect 56876 42764 56928 42770
rect 56876 42706 56928 42712
rect 56980 42362 57008 43182
rect 56968 42356 57020 42362
rect 56968 42298 57020 42304
rect 57336 42152 57388 42158
rect 57336 42094 57388 42100
rect 57244 41608 57296 41614
rect 57244 41550 57296 41556
rect 57152 41540 57204 41546
rect 57152 41482 57204 41488
rect 56784 41472 56836 41478
rect 56784 41414 56836 41420
rect 56796 41206 56824 41414
rect 57164 41206 57192 41482
rect 56784 41200 56836 41206
rect 56784 41142 56836 41148
rect 57152 41200 57204 41206
rect 57152 41142 57204 41148
rect 56796 39642 56824 41142
rect 56784 39636 56836 39642
rect 56784 39578 56836 39584
rect 56784 38208 56836 38214
rect 56784 38150 56836 38156
rect 56796 37874 56824 38150
rect 56784 37868 56836 37874
rect 56784 37810 56836 37816
rect 56796 37126 56824 37810
rect 57164 37806 57192 41142
rect 57256 41138 57284 41550
rect 57348 41274 57376 42094
rect 57336 41268 57388 41274
rect 57336 41210 57388 41216
rect 57244 41132 57296 41138
rect 57244 41074 57296 41080
rect 57256 40934 57284 41074
rect 57244 40928 57296 40934
rect 57244 40870 57296 40876
rect 57256 40730 57284 40870
rect 57244 40724 57296 40730
rect 57244 40666 57296 40672
rect 57336 39296 57388 39302
rect 57336 39238 57388 39244
rect 57348 38282 57376 39238
rect 57336 38276 57388 38282
rect 57336 38218 57388 38224
rect 56876 37800 56928 37806
rect 56876 37742 56928 37748
rect 57152 37800 57204 37806
rect 57152 37742 57204 37748
rect 56784 37120 56836 37126
rect 56784 37062 56836 37068
rect 56796 35766 56824 37062
rect 56888 36922 56916 37742
rect 57152 37188 57204 37194
rect 57152 37130 57204 37136
rect 56876 36916 56928 36922
rect 56876 36858 56928 36864
rect 57164 36582 57192 37130
rect 57244 36780 57296 36786
rect 57244 36722 57296 36728
rect 57152 36576 57204 36582
rect 57152 36518 57204 36524
rect 57060 36236 57112 36242
rect 57060 36178 57112 36184
rect 56968 36100 57020 36106
rect 56968 36042 57020 36048
rect 56784 35760 56836 35766
rect 56784 35702 56836 35708
rect 56980 35086 57008 36042
rect 57072 35086 57100 36178
rect 57164 35290 57192 36518
rect 57256 36378 57284 36722
rect 57336 36644 57388 36650
rect 57336 36586 57388 36592
rect 57244 36372 57296 36378
rect 57244 36314 57296 36320
rect 57152 35284 57204 35290
rect 57152 35226 57204 35232
rect 56968 35080 57020 35086
rect 56968 35022 57020 35028
rect 57060 35080 57112 35086
rect 57060 35022 57112 35028
rect 56692 34604 56744 34610
rect 56692 34546 56744 34552
rect 56968 34400 57020 34406
rect 56968 34342 57020 34348
rect 56980 34066 57008 34342
rect 56968 34060 57020 34066
rect 56968 34002 57020 34008
rect 56600 33516 56652 33522
rect 56600 33458 56652 33464
rect 56876 33516 56928 33522
rect 56876 33458 56928 33464
rect 56612 32842 56640 33458
rect 56600 32836 56652 32842
rect 56600 32778 56652 32784
rect 56508 32564 56560 32570
rect 56508 32506 56560 32512
rect 56612 32366 56640 32778
rect 56600 32360 56652 32366
rect 56600 32302 56652 32308
rect 56048 31952 56100 31958
rect 56048 31894 56100 31900
rect 56060 31346 56088 31894
rect 56612 31482 56640 32302
rect 56140 31476 56192 31482
rect 56140 31418 56192 31424
rect 56600 31476 56652 31482
rect 56600 31418 56652 31424
rect 56048 31340 56100 31346
rect 56048 31282 56100 31288
rect 56060 30938 56088 31282
rect 56152 31210 56180 31418
rect 56140 31204 56192 31210
rect 56140 31146 56192 31152
rect 56048 30932 56100 30938
rect 56048 30874 56100 30880
rect 56152 29646 56180 31146
rect 56324 31136 56376 31142
rect 56324 31078 56376 31084
rect 56336 30802 56364 31078
rect 56324 30796 56376 30802
rect 56324 30738 56376 30744
rect 56692 30252 56744 30258
rect 56692 30194 56744 30200
rect 56508 30048 56560 30054
rect 56508 29990 56560 29996
rect 56520 29714 56548 29990
rect 56508 29708 56560 29714
rect 56508 29650 56560 29656
rect 56140 29640 56192 29646
rect 56140 29582 56192 29588
rect 56324 29640 56376 29646
rect 56324 29582 56376 29588
rect 56336 29073 56364 29582
rect 56322 29064 56378 29073
rect 56322 28999 56378 29008
rect 56324 28552 56376 28558
rect 56324 28494 56376 28500
rect 56336 28082 56364 28494
rect 56324 28076 56376 28082
rect 56324 28018 56376 28024
rect 55956 27124 56008 27130
rect 55956 27066 56008 27072
rect 56600 26988 56652 26994
rect 56600 26930 56652 26936
rect 56508 25696 56560 25702
rect 56508 25638 56560 25644
rect 56520 25362 56548 25638
rect 56508 25356 56560 25362
rect 56508 25298 56560 25304
rect 56612 24818 56640 26930
rect 56600 24812 56652 24818
rect 56600 24754 56652 24760
rect 56508 24608 56560 24614
rect 56508 24550 56560 24556
rect 56520 24274 56548 24550
rect 56508 24268 56560 24274
rect 56508 24210 56560 24216
rect 56600 22432 56652 22438
rect 56600 22374 56652 22380
rect 56612 22098 56640 22374
rect 56600 22092 56652 22098
rect 56600 22034 56652 22040
rect 56324 16992 56376 16998
rect 56324 16934 56376 16940
rect 56336 16658 56364 16934
rect 56324 16652 56376 16658
rect 56324 16594 56376 16600
rect 56324 15904 56376 15910
rect 56324 15846 56376 15852
rect 56336 15570 56364 15846
rect 56324 15564 56376 15570
rect 56324 15506 56376 15512
rect 55680 15020 55732 15026
rect 55680 14962 55732 14968
rect 56324 14816 56376 14822
rect 56324 14758 56376 14764
rect 56336 14482 56364 14758
rect 56324 14476 56376 14482
rect 56324 14418 56376 14424
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 56704 10198 56732 30194
rect 56784 27464 56836 27470
rect 56784 27406 56836 27412
rect 56692 10192 56744 10198
rect 56692 10134 56744 10140
rect 56704 10062 56732 10134
rect 56692 10056 56744 10062
rect 56692 9998 56744 10004
rect 56692 9920 56744 9926
rect 56692 9862 56744 9868
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 56324 9376 56376 9382
rect 56324 9318 56376 9324
rect 56336 9042 56364 9318
rect 56704 9042 56732 9862
rect 56324 9036 56376 9042
rect 56324 8978 56376 8984
rect 56692 9036 56744 9042
rect 56692 8978 56744 8984
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 56324 6724 56376 6730
rect 56324 6666 56376 6672
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 56336 5778 56364 6666
rect 56600 6112 56652 6118
rect 56600 6054 56652 6060
rect 56324 5772 56376 5778
rect 56324 5714 56376 5720
rect 55496 5704 55548 5710
rect 55496 5646 55548 5652
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 55508 5234 55536 5646
rect 55496 5228 55548 5234
rect 55496 5170 55548 5176
rect 56324 5024 56376 5030
rect 56324 4966 56376 4972
rect 56336 4690 56364 4966
rect 56324 4684 56376 4690
rect 56324 4626 56376 4632
rect 56508 4684 56560 4690
rect 56508 4626 56560 4632
rect 55036 4616 55088 4622
rect 55036 4558 55088 4564
rect 55496 4616 55548 4622
rect 55496 4558 55548 4564
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 49976 4140 50028 4146
rect 49976 4082 50028 4088
rect 53840 4140 53892 4146
rect 53840 4082 53892 4088
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 48240 3058 48268 3470
rect 48320 3392 48372 3398
rect 48320 3334 48372 3340
rect 47584 3052 47636 3058
rect 47584 2994 47636 3000
rect 48228 3052 48280 3058
rect 48228 2994 48280 3000
rect 48332 800 48360 3334
rect 49988 3194 50016 4082
rect 50344 3936 50396 3942
rect 50344 3878 50396 3884
rect 53104 3936 53156 3942
rect 53104 3878 53156 3884
rect 50356 3602 50384 3878
rect 53116 3602 53144 3878
rect 50344 3596 50396 3602
rect 50344 3538 50396 3544
rect 50620 3596 50672 3602
rect 50620 3538 50672 3544
rect 53104 3596 53156 3602
rect 53104 3538 53156 3544
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 49976 3188 50028 3194
rect 49976 3130 50028 3136
rect 49608 2984 49660 2990
rect 49608 2926 49660 2932
rect 49620 800 49648 2926
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50632 1714 50660 3538
rect 52920 3528 52972 3534
rect 52920 3470 52972 3476
rect 52932 3058 52960 3470
rect 52920 3052 52972 3058
rect 52920 2994 52972 3000
rect 53852 2514 53880 4082
rect 54116 3596 54168 3602
rect 54116 3538 54168 3544
rect 54024 2984 54076 2990
rect 54024 2926 54076 2932
rect 54036 2650 54064 2926
rect 54024 2644 54076 2650
rect 54024 2586 54076 2592
rect 53840 2508 53892 2514
rect 53840 2450 53892 2456
rect 50264 1686 50660 1714
rect 50264 800 50292 1686
rect 54128 800 54156 3538
rect 54208 3392 54260 3398
rect 54208 3334 54260 3340
rect 54220 3126 54248 3334
rect 54208 3120 54260 3126
rect 54208 3062 54260 3068
rect 54760 2984 54812 2990
rect 54760 2926 54812 2932
rect 54772 800 54800 2926
rect 55048 2514 55076 4558
rect 55508 4146 55536 4558
rect 55496 4140 55548 4146
rect 55496 4082 55548 4088
rect 55404 3936 55456 3942
rect 55404 3878 55456 3884
rect 55036 2508 55088 2514
rect 55036 2450 55088 2456
rect 55416 2378 55444 3878
rect 56048 3460 56100 3466
rect 56048 3402 56100 3408
rect 55404 2372 55456 2378
rect 55404 2314 55456 2320
rect 56060 800 56088 3402
rect -10 0 102 800
rect 634 0 746 800
rect 1922 0 2034 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 21886 0 21998 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 25106 0 25218 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32834 0 32946 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 40562 0 40674 800
rect 41850 0 41962 800
rect 42494 0 42606 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 46358 0 46470 800
rect 47002 0 47114 800
rect 48290 0 48402 800
rect 49578 0 49690 800
rect 50222 0 50334 800
rect 51510 0 51622 800
rect 52798 0 52910 800
rect 54086 0 54198 800
rect 54730 0 54842 800
rect 56018 0 56130 800
rect 56520 105 56548 4626
rect 56612 4214 56640 6054
rect 56600 4208 56652 4214
rect 56600 4150 56652 4156
rect 56796 3738 56824 27406
rect 56888 18170 56916 33458
rect 56968 33312 57020 33318
rect 56968 33254 57020 33260
rect 56980 32434 57008 33254
rect 57072 32570 57100 35022
rect 57152 33312 57204 33318
rect 57152 33254 57204 33260
rect 57244 33312 57296 33318
rect 57244 33254 57296 33260
rect 57164 32978 57192 33254
rect 57256 33046 57284 33254
rect 57244 33040 57296 33046
rect 57244 32982 57296 32988
rect 57152 32972 57204 32978
rect 57152 32914 57204 32920
rect 57152 32768 57204 32774
rect 57152 32710 57204 32716
rect 57060 32564 57112 32570
rect 57060 32506 57112 32512
rect 57164 32434 57192 32710
rect 56968 32428 57020 32434
rect 56968 32370 57020 32376
rect 57152 32428 57204 32434
rect 57152 32370 57204 32376
rect 57348 30258 57376 36586
rect 57336 30252 57388 30258
rect 57336 30194 57388 30200
rect 56968 28484 57020 28490
rect 56968 28426 57020 28432
rect 56980 27606 57008 28426
rect 56968 27600 57020 27606
rect 56968 27542 57020 27548
rect 56968 26784 57020 26790
rect 56968 26726 57020 26732
rect 56980 26450 57008 26726
rect 56968 26444 57020 26450
rect 56968 26386 57020 26392
rect 57060 26308 57112 26314
rect 57060 26250 57112 26256
rect 57072 26042 57100 26250
rect 57060 26036 57112 26042
rect 57060 25978 57112 25984
rect 57440 25906 57468 45902
rect 57428 25900 57480 25906
rect 57428 25842 57480 25848
rect 57428 24812 57480 24818
rect 57428 24754 57480 24760
rect 57244 22432 57296 22438
rect 57244 22374 57296 22380
rect 57336 22432 57388 22438
rect 57336 22374 57388 22380
rect 57060 21344 57112 21350
rect 57060 21286 57112 21292
rect 57152 21344 57204 21350
rect 57152 21286 57204 21292
rect 57072 19922 57100 21286
rect 57164 19990 57192 21286
rect 57256 20874 57284 22374
rect 57348 22166 57376 22374
rect 57336 22160 57388 22166
rect 57336 22102 57388 22108
rect 57440 22094 57468 24754
rect 57532 22710 57560 51342
rect 57612 49156 57664 49162
rect 57612 49098 57664 49104
rect 57624 36650 57652 49098
rect 57716 43353 57744 57394
rect 57992 56914 58020 59200
rect 57980 56908 58032 56914
rect 57980 56850 58032 56856
rect 57980 56772 58032 56778
rect 57980 56714 58032 56720
rect 57992 55418 58020 56714
rect 57980 55412 58032 55418
rect 57980 55354 58032 55360
rect 58162 55176 58218 55185
rect 58162 55111 58218 55120
rect 58176 54738 58204 55111
rect 58164 54732 58216 54738
rect 58164 54674 58216 54680
rect 58162 53816 58218 53825
rect 58162 53751 58218 53760
rect 58176 53650 58204 53751
rect 58164 53644 58216 53650
rect 58164 53586 58216 53592
rect 57796 51400 57848 51406
rect 57796 51342 57848 51348
rect 57808 50454 57836 51342
rect 57886 51096 57942 51105
rect 57886 51031 57942 51040
rect 57796 50448 57848 50454
rect 57796 50390 57848 50396
rect 57900 50386 57928 51031
rect 57888 50380 57940 50386
rect 57888 50322 57940 50328
rect 57886 49056 57942 49065
rect 57886 48991 57942 49000
rect 57900 48210 57928 48991
rect 57888 48204 57940 48210
rect 57888 48146 57940 48152
rect 58072 47116 58124 47122
rect 58072 47058 58124 47064
rect 58084 46578 58112 47058
rect 58162 47016 58218 47025
rect 58162 46951 58164 46960
rect 58216 46951 58218 46960
rect 58164 46922 58216 46928
rect 58072 46572 58124 46578
rect 58072 46514 58124 46520
rect 57796 45960 57848 45966
rect 57796 45902 57848 45908
rect 57808 45014 57836 45902
rect 57886 45656 57942 45665
rect 57886 45591 57942 45600
rect 57796 45008 57848 45014
rect 57796 44950 57848 44956
rect 57900 44946 57928 45591
rect 57888 44940 57940 44946
rect 57888 44882 57940 44888
rect 57886 44296 57942 44305
rect 57886 44231 57942 44240
rect 57900 43858 57928 44231
rect 57888 43852 57940 43858
rect 57888 43794 57940 43800
rect 57702 43344 57758 43353
rect 57702 43279 57704 43288
rect 57756 43279 57758 43288
rect 57704 43250 57756 43256
rect 57612 36644 57664 36650
rect 57612 36586 57664 36592
rect 57716 36530 57744 43250
rect 57886 42936 57942 42945
rect 57886 42871 57942 42880
rect 57900 42770 57928 42871
rect 57888 42764 57940 42770
rect 57888 42706 57940 42712
rect 58072 42628 58124 42634
rect 58072 42570 58124 42576
rect 58084 42226 58112 42570
rect 58072 42220 58124 42226
rect 58072 42162 58124 42168
rect 57888 40044 57940 40050
rect 57888 39986 57940 39992
rect 57900 39545 57928 39986
rect 57886 39536 57942 39545
rect 57886 39471 57942 39480
rect 57796 39432 57848 39438
rect 57796 39374 57848 39380
rect 57624 36502 57744 36530
rect 57624 30258 57652 36502
rect 57808 35578 57836 39374
rect 57886 38856 57942 38865
rect 57886 38791 57942 38800
rect 57900 38418 57928 38791
rect 57888 38412 57940 38418
rect 57888 38354 57940 38360
rect 57980 37256 58032 37262
rect 57980 37198 58032 37204
rect 57992 36922 58020 37198
rect 57980 36916 58032 36922
rect 57980 36858 58032 36864
rect 57716 35550 57836 35578
rect 57612 30252 57664 30258
rect 57612 30194 57664 30200
rect 57520 22704 57572 22710
rect 57520 22646 57572 22652
rect 57624 22642 57652 30194
rect 57612 22636 57664 22642
rect 57612 22578 57664 22584
rect 57440 22066 57652 22094
rect 57244 20868 57296 20874
rect 57244 20810 57296 20816
rect 57152 19984 57204 19990
rect 57152 19926 57204 19932
rect 57060 19916 57112 19922
rect 57060 19858 57112 19864
rect 56888 18142 57008 18170
rect 56876 18080 56928 18086
rect 56876 18022 56928 18028
rect 56888 17746 56916 18022
rect 56876 17740 56928 17746
rect 56876 17682 56928 17688
rect 56980 16574 57008 18142
rect 57152 17604 57204 17610
rect 57152 17546 57204 17552
rect 57164 17338 57192 17546
rect 57152 17332 57204 17338
rect 57152 17274 57204 17280
rect 57060 17196 57112 17202
rect 57060 17138 57112 17144
rect 56888 16546 57008 16574
rect 56888 6798 56916 16546
rect 57072 16114 57100 17138
rect 57152 16516 57204 16522
rect 57152 16458 57204 16464
rect 57164 16250 57192 16458
rect 57152 16244 57204 16250
rect 57152 16186 57204 16192
rect 57060 16108 57112 16114
rect 57060 16050 57112 16056
rect 56968 15428 57020 15434
rect 56968 15370 57020 15376
rect 56980 15162 57008 15370
rect 57072 15366 57100 16050
rect 57060 15360 57112 15366
rect 57060 15302 57112 15308
rect 56968 15156 57020 15162
rect 56968 15098 57020 15104
rect 57336 15020 57388 15026
rect 57336 14962 57388 14968
rect 56968 14340 57020 14346
rect 56968 14282 57020 14288
rect 56980 14074 57008 14282
rect 56968 14068 57020 14074
rect 56968 14010 57020 14016
rect 57152 13932 57204 13938
rect 57152 13874 57204 13880
rect 56876 6792 56928 6798
rect 56876 6734 56928 6740
rect 57060 6656 57112 6662
rect 57060 6598 57112 6604
rect 57072 5302 57100 6598
rect 57060 5296 57112 5302
rect 57060 5238 57112 5244
rect 57164 3942 57192 13874
rect 57244 9988 57296 9994
rect 57244 9930 57296 9936
rect 57256 9625 57284 9930
rect 57242 9616 57298 9625
rect 57242 9551 57298 9560
rect 57348 6118 57376 14962
rect 57336 6112 57388 6118
rect 57336 6054 57388 6060
rect 57152 3936 57204 3942
rect 57152 3878 57204 3884
rect 56784 3732 56836 3738
rect 56784 3674 56836 3680
rect 56796 3058 56824 3674
rect 57624 3670 57652 22066
rect 57716 21554 57744 35550
rect 57886 34776 57942 34785
rect 57886 34711 57942 34720
rect 57794 34096 57850 34105
rect 57900 34066 57928 34711
rect 58072 34400 58124 34406
rect 58072 34342 58124 34348
rect 58084 34134 58112 34342
rect 58072 34128 58124 34134
rect 58072 34070 58124 34076
rect 57794 34031 57850 34040
rect 57888 34060 57940 34066
rect 57808 32978 57836 34031
rect 57888 34002 57940 34008
rect 57796 32972 57848 32978
rect 57796 32914 57848 32920
rect 57794 32736 57850 32745
rect 57794 32671 57850 32680
rect 57808 28626 57836 32671
rect 57886 31376 57942 31385
rect 57886 31311 57942 31320
rect 57900 29714 57928 31311
rect 58162 30696 58218 30705
rect 57980 30660 58032 30666
rect 58162 30631 58164 30640
rect 57980 30602 58032 30608
rect 58216 30631 58218 30640
rect 58164 30602 58216 30608
rect 57992 30326 58020 30602
rect 57980 30320 58032 30326
rect 57980 30262 58032 30268
rect 57888 29708 57940 29714
rect 57888 29650 57940 29656
rect 57796 28620 57848 28626
rect 57796 28562 57848 28568
rect 58162 26616 58218 26625
rect 58162 26551 58218 26560
rect 58176 26450 58204 26551
rect 58164 26444 58216 26450
rect 58164 26386 58216 26392
rect 58162 25936 58218 25945
rect 58162 25871 58218 25880
rect 58072 25696 58124 25702
rect 58072 25638 58124 25644
rect 58084 25430 58112 25638
rect 58072 25424 58124 25430
rect 58072 25366 58124 25372
rect 58176 25362 58204 25871
rect 58164 25356 58216 25362
rect 58164 25298 58216 25304
rect 58072 24608 58124 24614
rect 58072 24550 58124 24556
rect 58162 24576 58218 24585
rect 58084 24342 58112 24550
rect 58162 24511 58218 24520
rect 58072 24336 58124 24342
rect 58072 24278 58124 24284
rect 58176 24274 58204 24511
rect 58164 24268 58216 24274
rect 58164 24210 58216 24216
rect 57886 22536 57942 22545
rect 57886 22471 57942 22480
rect 57900 22098 57928 22471
rect 57888 22092 57940 22098
rect 57888 22034 57940 22040
rect 57704 21548 57756 21554
rect 57704 21490 57756 21496
rect 57794 21176 57850 21185
rect 57794 21111 57850 21120
rect 57808 19922 57836 21111
rect 57888 21004 57940 21010
rect 57888 20946 57940 20952
rect 57796 19916 57848 19922
rect 57796 19858 57848 19864
rect 57900 19825 57928 20946
rect 58072 20936 58124 20942
rect 58072 20878 58124 20884
rect 58084 20466 58112 20878
rect 58072 20460 58124 20466
rect 58072 20402 58124 20408
rect 57886 19816 57942 19825
rect 57886 19751 57942 19760
rect 58162 17776 58218 17785
rect 58162 17711 58164 17720
rect 58216 17711 58218 17720
rect 58164 17682 58216 17688
rect 57796 16652 57848 16658
rect 57796 16594 57848 16600
rect 57808 16425 57836 16594
rect 57794 16416 57850 16425
rect 57794 16351 57850 16360
rect 57888 15564 57940 15570
rect 57888 15506 57940 15512
rect 57796 15360 57848 15366
rect 57796 15302 57848 15308
rect 57808 4146 57836 15302
rect 57900 15065 57928 15506
rect 57886 15056 57942 15065
rect 57886 14991 57942 15000
rect 58162 14376 58218 14385
rect 58162 14311 58164 14320
rect 58216 14311 58218 14320
rect 58164 14282 58216 14288
rect 57888 9036 57940 9042
rect 57888 8978 57940 8984
rect 57900 8265 57928 8978
rect 57886 8256 57942 8265
rect 57886 8191 57942 8200
rect 58162 6216 58218 6225
rect 58162 6151 58218 6160
rect 57980 6112 58032 6118
rect 57980 6054 58032 6060
rect 57992 5778 58020 6054
rect 58176 5778 58204 6151
rect 57980 5772 58032 5778
rect 57980 5714 58032 5720
rect 58164 5772 58216 5778
rect 58164 5714 58216 5720
rect 58624 5160 58676 5166
rect 58624 5102 58676 5108
rect 57980 4548 58032 4554
rect 57980 4490 58032 4496
rect 57796 4140 57848 4146
rect 57796 4082 57848 4088
rect 57704 4072 57756 4078
rect 57704 4014 57756 4020
rect 57612 3664 57664 3670
rect 57612 3606 57664 3612
rect 56968 3460 57020 3466
rect 56968 3402 57020 3408
rect 56980 3194 57008 3402
rect 56968 3188 57020 3194
rect 56968 3130 57020 3136
rect 56784 3052 56836 3058
rect 56784 2994 56836 3000
rect 57336 2372 57388 2378
rect 57336 2314 57388 2320
rect 57348 800 57376 2314
rect 57716 2145 57744 4014
rect 57888 3596 57940 3602
rect 57888 3538 57940 3544
rect 57702 2136 57758 2145
rect 57702 2071 57758 2080
rect 57900 1465 57928 3538
rect 57992 3194 58020 4490
rect 58072 3528 58124 3534
rect 58072 3470 58124 3476
rect 57980 3188 58032 3194
rect 57980 3130 58032 3136
rect 58084 2650 58112 3470
rect 58072 2644 58124 2650
rect 58072 2586 58124 2592
rect 57886 1456 57942 1465
rect 57886 1391 57942 1400
rect 58636 800 58664 5102
rect 56506 96 56562 105
rect 56506 31 56562 40
rect 57306 0 57418 800
rect 58594 0 58706 800
rect 59238 0 59350 800
<< via2 >>
rect 1490 55800 1546 55856
rect 2778 57840 2834 57896
rect 3974 57160 4030 57216
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 2778 54440 2834 54496
rect 3238 52400 3294 52456
rect 2962 49000 3018 49056
rect 3422 49716 3424 49736
rect 3424 49716 3476 49736
rect 3476 49716 3478 49736
rect 3422 49680 3478 49716
rect 2778 39480 2834 39536
rect 2778 29960 2834 30016
rect 2778 26560 2834 26616
rect 2778 24520 2834 24576
rect 2778 21800 2834 21856
rect 2778 20440 2834 20496
rect 2778 18400 2834 18456
rect 2778 17076 2780 17096
rect 2780 17076 2832 17096
rect 2832 17076 2834 17096
rect 2778 17040 2834 17076
rect 2778 13640 2834 13696
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 2778 8200 2834 8256
rect 2778 6840 2834 6896
rect 3422 28600 3478 28656
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3974 12280 4030 12336
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3422 8880 3478 8936
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2778 4120 2834 4176
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3238 5480 3294 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 2870 3440 2926 3496
rect 2778 2080 2834 2136
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 20442 41656 20498 41712
rect 20810 41556 20812 41576
rect 20812 41556 20864 41576
rect 20864 41556 20866 41576
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 20810 41520 20866 41556
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 21914 41556 21916 41576
rect 21916 41556 21968 41576
rect 21968 41556 21970 41576
rect 21914 41520 21970 41556
rect 22558 41656 22614 41712
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 28906 43288 28962 43344
rect 29550 27512 29606 27568
rect 30194 26308 30250 26344
rect 30194 26288 30196 26308
rect 30196 26288 30248 26308
rect 30248 26288 30250 26308
rect 31206 41792 31262 41848
rect 30930 38256 30986 38312
rect 31114 38664 31170 38720
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 31298 38664 31354 38720
rect 31298 38256 31354 38312
rect 31022 36760 31078 36816
rect 30746 26324 30748 26344
rect 30748 26324 30800 26344
rect 30800 26324 30802 26344
rect 30746 26288 30802 26324
rect 30930 26324 30932 26344
rect 30932 26324 30984 26344
rect 30984 26324 30986 26344
rect 30930 26288 30986 26324
rect 33506 47116 33562 47152
rect 33506 47096 33508 47116
rect 33508 47096 33560 47116
rect 33560 47096 33562 47116
rect 34150 41792 34206 41848
rect 33414 38800 33470 38856
rect 33598 38664 33654 38720
rect 34242 38820 34298 38856
rect 34242 38800 34244 38820
rect 34244 38800 34296 38820
rect 34296 38800 34298 38820
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 42614 55392 42670 55448
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34610 38664 34666 38720
rect 34518 38392 34574 38448
rect 34334 38256 34390 38312
rect 34518 38256 34574 38312
rect 31574 27784 31630 27840
rect 32126 27820 32128 27840
rect 32128 27820 32180 27840
rect 32180 27820 32182 27840
rect 32126 27784 32182 27820
rect 31850 26324 31852 26344
rect 31852 26324 31904 26344
rect 31904 26324 31906 26344
rect 31850 26288 31906 26324
rect 33690 29572 33746 29608
rect 33690 29552 33692 29572
rect 33692 29552 33744 29572
rect 33744 29552 33746 29572
rect 33506 29028 33562 29064
rect 33506 29008 33508 29028
rect 33508 29008 33560 29028
rect 33560 29008 33562 29028
rect 32862 27548 32864 27568
rect 32864 27548 32916 27568
rect 32916 27548 32918 27568
rect 32862 27512 32918 27548
rect 34058 28192 34114 28248
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 35990 44396 36046 44432
rect 35990 44376 35992 44396
rect 35992 44376 36044 44396
rect 36044 44376 36046 44396
rect 36450 45328 36506 45384
rect 36450 45228 36452 45248
rect 36452 45228 36504 45248
rect 36504 45228 36506 45248
rect 36450 45192 36506 45228
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 35346 38612 35402 38668
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35162 38412 35218 38448
rect 35162 38392 35164 38412
rect 35164 38392 35216 38412
rect 35216 38392 35218 38412
rect 35346 38256 35402 38312
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 36542 36780 36598 36816
rect 36542 36760 36544 36780
rect 36544 36760 36596 36780
rect 36596 36760 36598 36780
rect 36082 33904 36138 33960
rect 39670 46996 39672 47016
rect 39672 46996 39724 47016
rect 39724 46996 39726 47016
rect 39670 46960 39726 46996
rect 39210 46572 39266 46608
rect 39210 46552 39212 46572
rect 39212 46552 39264 46572
rect 39264 46552 39266 46572
rect 37922 45348 37978 45384
rect 37922 45328 37924 45348
rect 37924 45328 37976 45348
rect 37976 45328 37978 45348
rect 38198 45228 38200 45248
rect 38200 45228 38252 45248
rect 38252 45228 38254 45248
rect 38198 45192 38254 45228
rect 37094 38800 37150 38856
rect 37370 36780 37426 36816
rect 37370 36760 37372 36780
rect 37372 36760 37424 36780
rect 37424 36760 37426 36780
rect 37186 33496 37242 33552
rect 39946 45500 39948 45520
rect 39948 45500 40000 45520
rect 40000 45500 40002 45520
rect 39946 45464 40002 45500
rect 39026 43868 39028 43888
rect 39028 43868 39080 43888
rect 39080 43868 39082 43888
rect 39026 43832 39082 43868
rect 38382 37712 38438 37768
rect 39394 38972 39396 38992
rect 39396 38972 39448 38992
rect 39448 38972 39450 38992
rect 39394 38936 39450 38972
rect 39394 38820 39450 38856
rect 39394 38800 39396 38820
rect 39396 38800 39448 38820
rect 39448 38800 39450 38820
rect 40314 43560 40370 43616
rect 39578 38004 39634 38040
rect 39578 37984 39580 38004
rect 39580 37984 39632 38004
rect 39632 37984 39634 38004
rect 40866 46960 40922 47016
rect 40682 43968 40738 44024
rect 40958 44648 41014 44704
rect 41050 44240 41106 44296
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 56506 58520 56562 58576
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 41510 46552 41566 46608
rect 41970 46980 42026 47016
rect 41970 46960 41972 46980
rect 41972 46960 42024 46980
rect 42024 46960 42026 46980
rect 40590 38800 40646 38856
rect 40682 37712 40738 37768
rect 40406 34448 40462 34504
rect 39578 25916 39580 25936
rect 39580 25916 39632 25936
rect 39632 25916 39634 25936
rect 39578 25880 39634 25916
rect 40682 34448 40738 34504
rect 41602 42608 41658 42664
rect 42154 43188 42156 43208
rect 42156 43188 42208 43208
rect 42208 43188 42210 43208
rect 42154 43152 42210 43188
rect 41326 38936 41382 38992
rect 42430 44648 42486 44704
rect 42982 43832 43038 43888
rect 42982 43424 43038 43480
rect 41786 38528 41842 38584
rect 42522 35148 42578 35184
rect 42522 35128 42524 35148
rect 42524 35128 42576 35148
rect 42576 35128 42578 35148
rect 42798 37868 42854 37904
rect 42798 37848 42800 37868
rect 42800 37848 42852 37868
rect 42852 37848 42854 37868
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 45374 46996 45376 47016
rect 45376 46996 45428 47016
rect 45428 46996 45430 47016
rect 45374 46960 45430 46996
rect 43626 43424 43682 43480
rect 44086 43152 44142 43208
rect 42798 34620 42800 34640
rect 42800 34620 42852 34640
rect 42852 34620 42854 34640
rect 42798 34584 42854 34620
rect 40682 28328 40738 28384
rect 40590 27376 40646 27432
rect 40314 25916 40316 25936
rect 40316 25916 40368 25936
rect 40368 25916 40370 25936
rect 40314 25880 40370 25916
rect 42706 29552 42762 29608
rect 43902 33260 43904 33280
rect 43904 33260 43956 33280
rect 43956 33260 43958 33280
rect 43902 33224 43958 33260
rect 44270 35128 44326 35184
rect 44178 34604 44234 34640
rect 44178 34584 44180 34604
rect 44180 34584 44232 34604
rect 44232 34584 44234 34604
rect 43718 29572 43774 29608
rect 43718 29552 43720 29572
rect 43720 29552 43772 29572
rect 43772 29552 43774 29572
rect 42338 27412 42340 27432
rect 42340 27412 42392 27432
rect 42392 27412 42394 27432
rect 42338 27376 42394 27412
rect 40682 24792 40738 24848
rect 43626 24676 43682 24712
rect 43626 24656 43628 24676
rect 43628 24656 43680 24676
rect 43680 24656 43682 24676
rect 45834 47504 45890 47560
rect 44638 43444 44694 43480
rect 44638 43424 44640 43444
rect 44640 43424 44692 43444
rect 44692 43424 44694 43444
rect 45190 44104 45246 44160
rect 45006 42644 45008 42664
rect 45008 42644 45060 42664
rect 45060 42644 45062 42664
rect 45006 42608 45062 42644
rect 45650 43852 45706 43888
rect 45834 44260 45890 44296
rect 45834 44240 45836 44260
rect 45836 44240 45888 44260
rect 45888 44240 45890 44260
rect 45650 43832 45652 43852
rect 45652 43832 45704 43852
rect 45704 43832 45706 43852
rect 46018 43560 46074 43616
rect 46662 44240 46718 44296
rect 46570 44104 46626 44160
rect 45282 37984 45338 38040
rect 46386 38528 46442 38584
rect 45742 34448 45798 34504
rect 47858 47504 47914 47560
rect 47582 43968 47638 44024
rect 47766 43832 47822 43888
rect 48134 45464 48190 45520
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 47674 37868 47730 37904
rect 47674 37848 47676 37868
rect 47676 37848 47728 37868
rect 47728 37848 47730 37868
rect 46386 24812 46442 24848
rect 46386 24792 46388 24812
rect 46388 24792 46440 24812
rect 46440 24792 46442 24812
rect 49422 44956 49424 44976
rect 49424 44956 49476 44976
rect 49476 44956 49478 44976
rect 49422 44920 49478 44956
rect 48318 39908 48374 39944
rect 48318 39888 48320 39908
rect 48320 39888 48372 39908
rect 48372 39888 48374 39908
rect 49698 44376 49754 44432
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 49054 33904 49110 33960
rect 49054 33224 49110 33280
rect 49238 33360 49294 33416
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 55494 44956 55496 44976
rect 55496 44956 55548 44976
rect 55548 44956 55550 44976
rect 55494 44920 55550 44956
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 49790 37984 49846 38040
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 49882 34992 49938 35048
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50250 34620 50252 34640
rect 50252 34620 50304 34640
rect 50304 34620 50306 34640
rect 50250 34584 50306 34620
rect 49974 33904 50030 33960
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 49974 32292 50030 32328
rect 49974 32272 49976 32292
rect 49976 32272 50028 32292
rect 50028 32272 50030 32292
rect 48042 28328 48098 28384
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 51446 34604 51502 34640
rect 51446 34584 51448 34604
rect 51448 34584 51500 34604
rect 51500 34584 51502 34604
rect 51722 34992 51778 35048
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 53930 39908 53986 39944
rect 53930 39888 53932 39908
rect 53932 39888 53984 39908
rect 53984 39888 53986 39908
rect 55218 27920 55274 27976
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 47950 24692 47952 24712
rect 47952 24692 48004 24712
rect 48004 24692 48006 24712
rect 47950 24656 48006 24692
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 57334 55800 57390 55856
rect 56322 29008 56378 29064
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 58162 55120 58218 55176
rect 58162 53760 58218 53816
rect 57886 51040 57942 51096
rect 57886 49000 57942 49056
rect 58162 46980 58218 47016
rect 58162 46960 58164 46980
rect 58164 46960 58216 46980
rect 58216 46960 58218 46980
rect 57886 45600 57942 45656
rect 57886 44240 57942 44296
rect 57702 43308 57758 43344
rect 57702 43288 57704 43308
rect 57704 43288 57756 43308
rect 57756 43288 57758 43308
rect 57886 42880 57942 42936
rect 57886 39480 57942 39536
rect 57886 38800 57942 38856
rect 57242 9560 57298 9616
rect 57886 34720 57942 34776
rect 57794 34040 57850 34096
rect 57794 32680 57850 32736
rect 57886 31320 57942 31376
rect 58162 30660 58218 30696
rect 58162 30640 58164 30660
rect 58164 30640 58216 30660
rect 58216 30640 58218 30660
rect 58162 26560 58218 26616
rect 58162 25880 58218 25936
rect 58162 24520 58218 24576
rect 57886 22480 57942 22536
rect 57794 21120 57850 21176
rect 57886 19760 57942 19816
rect 58162 17740 58218 17776
rect 58162 17720 58164 17740
rect 58164 17720 58216 17740
rect 58216 17720 58218 17740
rect 57794 16360 57850 16416
rect 57886 15000 57942 15056
rect 58162 14340 58218 14376
rect 58162 14320 58164 14340
rect 58164 14320 58216 14340
rect 58216 14320 58218 14340
rect 57886 8200 57942 8256
rect 58162 6160 58218 6216
rect 57702 2080 57758 2136
rect 57886 1400 57942 1456
rect 56506 40 56562 96
<< metal3 >>
rect 0 59108 800 59348
rect 56501 58578 56567 58581
rect 59200 58578 60000 58668
rect 56501 58576 60000 58578
rect 56501 58520 56506 58576
rect 56562 58520 60000 58576
rect 56501 58518 60000 58520
rect 56501 58515 56567 58518
rect 59200 58428 60000 58518
rect 0 57898 800 57988
rect 2773 57898 2839 57901
rect 0 57896 2839 57898
rect 0 57840 2778 57896
rect 2834 57840 2839 57896
rect 0 57838 2839 57840
rect 0 57748 800 57838
rect 2773 57835 2839 57838
rect 19568 57696 19888 57697
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 57631 19888 57632
rect 50288 57696 50608 57697
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 57631 50608 57632
rect 0 57218 800 57308
rect 3969 57218 4035 57221
rect 0 57216 4035 57218
rect 0 57160 3974 57216
rect 4030 57160 4035 57216
rect 0 57158 4035 57160
rect 0 57068 800 57158
rect 3969 57155 4035 57158
rect 4208 57152 4528 57153
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 57087 4528 57088
rect 34928 57152 35248 57153
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 57087 35248 57088
rect 59200 57068 60000 57308
rect 19568 56608 19888 56609
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 56543 19888 56544
rect 50288 56608 50608 56609
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 56543 50608 56544
rect 4208 56064 4528 56065
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 55999 4528 56000
rect 34928 56064 35248 56065
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 55999 35248 56000
rect 0 55858 800 55948
rect 1485 55858 1551 55861
rect 0 55856 1551 55858
rect 0 55800 1490 55856
rect 1546 55800 1551 55856
rect 0 55798 1551 55800
rect 0 55708 800 55798
rect 1485 55795 1551 55798
rect 57329 55858 57395 55861
rect 59200 55858 60000 55948
rect 57329 55856 60000 55858
rect 57329 55800 57334 55856
rect 57390 55800 60000 55856
rect 57329 55798 60000 55800
rect 57329 55795 57395 55798
rect 59200 55708 60000 55798
rect 19568 55520 19888 55521
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 55455 19888 55456
rect 50288 55520 50608 55521
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 55455 50608 55456
rect 42609 55452 42675 55453
rect 42558 55450 42564 55452
rect 42518 55390 42564 55450
rect 42628 55448 42675 55452
rect 42670 55392 42675 55448
rect 42558 55388 42564 55390
rect 42628 55388 42675 55392
rect 42609 55387 42675 55388
rect 58157 55178 58223 55181
rect 59200 55178 60000 55268
rect 58157 55176 60000 55178
rect 58157 55120 58162 55176
rect 58218 55120 60000 55176
rect 58157 55118 60000 55120
rect 58157 55115 58223 55118
rect 59200 55028 60000 55118
rect 4208 54976 4528 54977
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 54911 4528 54912
rect 34928 54976 35248 54977
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 54911 35248 54912
rect 0 54498 800 54588
rect 2773 54498 2839 54501
rect 0 54496 2839 54498
rect 0 54440 2778 54496
rect 2834 54440 2839 54496
rect 0 54438 2839 54440
rect 0 54348 800 54438
rect 2773 54435 2839 54438
rect 19568 54432 19888 54433
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 54367 19888 54368
rect 50288 54432 50608 54433
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 54367 50608 54368
rect 4208 53888 4528 53889
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 53823 4528 53824
rect 34928 53888 35248 53889
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 53823 35248 53824
rect 58157 53818 58223 53821
rect 59200 53818 60000 53908
rect 58157 53816 60000 53818
rect 58157 53760 58162 53816
rect 58218 53760 60000 53816
rect 58157 53758 60000 53760
rect 58157 53755 58223 53758
rect 59200 53668 60000 53758
rect 19568 53344 19888 53345
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 53279 19888 53280
rect 50288 53344 50608 53345
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 53279 50608 53280
rect 0 52988 800 53228
rect 4208 52800 4528 52801
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 52735 4528 52736
rect 34928 52800 35248 52801
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 52735 35248 52736
rect 0 52458 800 52548
rect 3233 52458 3299 52461
rect 0 52456 3299 52458
rect 0 52400 3238 52456
rect 3294 52400 3299 52456
rect 0 52398 3299 52400
rect 0 52308 800 52398
rect 3233 52395 3299 52398
rect 59200 52308 60000 52548
rect 19568 52256 19888 52257
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 52191 19888 52192
rect 50288 52256 50608 52257
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 52191 50608 52192
rect 4208 51712 4528 51713
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 51647 4528 51648
rect 34928 51712 35248 51713
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 51647 35248 51648
rect 0 50948 800 51188
rect 19568 51168 19888 51169
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 51103 19888 51104
rect 50288 51168 50608 51169
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 51103 50608 51104
rect 57881 51098 57947 51101
rect 59200 51098 60000 51188
rect 57881 51096 60000 51098
rect 57881 51040 57886 51096
rect 57942 51040 60000 51096
rect 57881 51038 60000 51040
rect 57881 51035 57947 51038
rect 59200 50948 60000 51038
rect 4208 50624 4528 50625
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 50559 4528 50560
rect 34928 50624 35248 50625
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 50559 35248 50560
rect 59200 50268 60000 50508
rect 19568 50080 19888 50081
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 50015 19888 50016
rect 50288 50080 50608 50081
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 50015 50608 50016
rect 0 49738 800 49828
rect 3417 49738 3483 49741
rect 0 49736 3483 49738
rect 0 49680 3422 49736
rect 3478 49680 3483 49736
rect 0 49678 3483 49680
rect 0 49588 800 49678
rect 3417 49675 3483 49678
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 0 49058 800 49148
rect 2957 49058 3023 49061
rect 0 49056 3023 49058
rect 0 49000 2962 49056
rect 3018 49000 3023 49056
rect 0 48998 3023 49000
rect 0 48908 800 48998
rect 2957 48995 3023 48998
rect 57881 49058 57947 49061
rect 59200 49058 60000 49148
rect 57881 49056 60000 49058
rect 57881 49000 57886 49056
rect 57942 49000 60000 49056
rect 57881 48998 60000 49000
rect 57881 48995 57947 48998
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 48927 19888 48928
rect 50288 48992 50608 48993
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 48927 50608 48928
rect 59200 48908 60000 48998
rect 4208 48448 4528 48449
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 50288 47904 50608 47905
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 47839 50608 47840
rect 0 47548 800 47788
rect 59200 47698 60000 47788
rect 41370 47638 60000 47698
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 33501 47154 33567 47157
rect 41370 47154 41430 47638
rect 45829 47562 45895 47565
rect 47853 47562 47919 47565
rect 45829 47560 47919 47562
rect 45829 47504 45834 47560
rect 45890 47504 47858 47560
rect 47914 47504 47919 47560
rect 59200 47548 60000 47638
rect 45829 47502 47919 47504
rect 45829 47499 45895 47502
rect 47853 47499 47919 47502
rect 33501 47152 41430 47154
rect 33501 47096 33506 47152
rect 33562 47096 41430 47152
rect 33501 47094 41430 47096
rect 33501 47091 33567 47094
rect 39665 47018 39731 47021
rect 40861 47018 40927 47021
rect 39665 47016 40927 47018
rect 39665 46960 39670 47016
rect 39726 46960 40866 47016
rect 40922 46960 40927 47016
rect 39665 46958 40927 46960
rect 39665 46955 39731 46958
rect 40861 46955 40927 46958
rect 41965 47018 42031 47021
rect 45369 47018 45435 47021
rect 41965 47016 45435 47018
rect 41965 46960 41970 47016
rect 42026 46960 45374 47016
rect 45430 46960 45435 47016
rect 41965 46958 45435 46960
rect 41965 46955 42031 46958
rect 45369 46955 45435 46958
rect 58157 47018 58223 47021
rect 59200 47018 60000 47108
rect 58157 47016 60000 47018
rect 58157 46960 58162 47016
rect 58218 46960 60000 47016
rect 58157 46958 60000 46960
rect 58157 46955 58223 46958
rect 59200 46868 60000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 50288 46816 50608 46817
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 46751 50608 46752
rect 39205 46610 39271 46613
rect 41505 46610 41571 46613
rect 39205 46608 41571 46610
rect 39205 46552 39210 46608
rect 39266 46552 41510 46608
rect 41566 46552 41571 46608
rect 39205 46550 41571 46552
rect 39205 46547 39271 46550
rect 41505 46547 41571 46550
rect 0 46188 800 46428
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 50288 45728 50608 45729
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 45663 50608 45664
rect 57881 45658 57947 45661
rect 59200 45658 60000 45748
rect 57881 45656 60000 45658
rect 57881 45600 57886 45656
rect 57942 45600 60000 45656
rect 57881 45598 60000 45600
rect 57881 45595 57947 45598
rect 39941 45522 40007 45525
rect 48129 45522 48195 45525
rect 39941 45520 48195 45522
rect 39941 45464 39946 45520
rect 40002 45464 48134 45520
rect 48190 45464 48195 45520
rect 59200 45508 60000 45598
rect 39941 45462 48195 45464
rect 39941 45459 40007 45462
rect 48129 45459 48195 45462
rect 36445 45386 36511 45389
rect 37917 45386 37983 45389
rect 36445 45384 37983 45386
rect 36445 45328 36450 45384
rect 36506 45328 37922 45384
rect 37978 45328 37983 45384
rect 36445 45326 37983 45328
rect 36445 45323 36511 45326
rect 37917 45323 37983 45326
rect 36445 45250 36511 45253
rect 38193 45250 38259 45253
rect 36445 45248 38259 45250
rect 36445 45192 36450 45248
rect 36506 45192 38198 45248
rect 38254 45192 38259 45248
rect 36445 45190 38259 45192
rect 36445 45187 36511 45190
rect 38193 45187 38259 45190
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44828 800 45068
rect 49417 44978 49483 44981
rect 55489 44978 55555 44981
rect 49417 44976 55555 44978
rect 49417 44920 49422 44976
rect 49478 44920 55494 44976
rect 55550 44920 55555 44976
rect 49417 44918 55555 44920
rect 49417 44915 49483 44918
rect 55489 44915 55555 44918
rect 40953 44706 41019 44709
rect 42425 44706 42491 44709
rect 40953 44704 42491 44706
rect 40953 44648 40958 44704
rect 41014 44648 42430 44704
rect 42486 44648 42491 44704
rect 40953 44646 42491 44648
rect 40953 44643 41019 44646
rect 42425 44643 42491 44646
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 50288 44640 50608 44641
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 44575 50608 44576
rect 35985 44434 36051 44437
rect 49693 44434 49759 44437
rect 35985 44432 49759 44434
rect 0 44148 800 44388
rect 35985 44376 35990 44432
rect 36046 44376 49698 44432
rect 49754 44376 49759 44432
rect 35985 44374 49759 44376
rect 35985 44371 36051 44374
rect 49693 44371 49759 44374
rect 41045 44298 41111 44301
rect 45829 44298 45895 44301
rect 46657 44298 46723 44301
rect 41045 44296 46723 44298
rect 41045 44240 41050 44296
rect 41106 44240 45834 44296
rect 45890 44240 46662 44296
rect 46718 44240 46723 44296
rect 41045 44238 46723 44240
rect 41045 44235 41111 44238
rect 45829 44235 45895 44238
rect 46657 44235 46723 44238
rect 57881 44298 57947 44301
rect 59200 44298 60000 44388
rect 57881 44296 60000 44298
rect 57881 44240 57886 44296
rect 57942 44240 60000 44296
rect 57881 44238 60000 44240
rect 57881 44235 57947 44238
rect 45185 44162 45251 44165
rect 46565 44162 46631 44165
rect 45185 44160 46631 44162
rect 45185 44104 45190 44160
rect 45246 44104 46570 44160
rect 46626 44104 46631 44160
rect 59200 44148 60000 44238
rect 45185 44102 46631 44104
rect 45185 44099 45251 44102
rect 46565 44099 46631 44102
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 40677 44026 40743 44029
rect 47577 44026 47643 44029
rect 40677 44024 47643 44026
rect 40677 43968 40682 44024
rect 40738 43968 47582 44024
rect 47638 43968 47643 44024
rect 40677 43966 47643 43968
rect 40677 43963 40743 43966
rect 47577 43963 47643 43966
rect 39021 43890 39087 43893
rect 42977 43890 43043 43893
rect 39021 43888 43043 43890
rect 39021 43832 39026 43888
rect 39082 43832 42982 43888
rect 43038 43832 43043 43888
rect 39021 43830 43043 43832
rect 39021 43827 39087 43830
rect 42977 43827 43043 43830
rect 45645 43890 45711 43893
rect 47761 43890 47827 43893
rect 45645 43888 47827 43890
rect 45645 43832 45650 43888
rect 45706 43832 47766 43888
rect 47822 43832 47827 43888
rect 45645 43830 47827 43832
rect 45645 43827 45711 43830
rect 47761 43827 47827 43830
rect 40309 43618 40375 43621
rect 46013 43618 46079 43621
rect 40309 43616 46079 43618
rect 40309 43560 40314 43616
rect 40370 43560 46018 43616
rect 46074 43560 46079 43616
rect 40309 43558 46079 43560
rect 40309 43555 40375 43558
rect 46013 43555 46079 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 50288 43552 50608 43553
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 43487 50608 43488
rect 42977 43482 43043 43485
rect 43621 43482 43687 43485
rect 44633 43482 44699 43485
rect 42977 43480 44699 43482
rect 42977 43424 42982 43480
rect 43038 43424 43626 43480
rect 43682 43424 44638 43480
rect 44694 43424 44699 43480
rect 42977 43422 44699 43424
rect 42977 43419 43043 43422
rect 43621 43419 43687 43422
rect 44633 43419 44699 43422
rect 28901 43346 28967 43349
rect 57697 43346 57763 43349
rect 28901 43344 57763 43346
rect 28901 43288 28906 43344
rect 28962 43288 57702 43344
rect 57758 43288 57763 43344
rect 28901 43286 57763 43288
rect 28901 43283 28967 43286
rect 57697 43283 57763 43286
rect 42149 43210 42215 43213
rect 44081 43210 44147 43213
rect 42149 43208 44147 43210
rect 42149 43152 42154 43208
rect 42210 43152 44086 43208
rect 44142 43152 44147 43208
rect 42149 43150 44147 43152
rect 42149 43147 42215 43150
rect 44081 43147 44147 43150
rect 0 42788 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 57881 42938 57947 42941
rect 59200 42938 60000 43028
rect 57881 42936 60000 42938
rect 57881 42880 57886 42936
rect 57942 42880 60000 42936
rect 57881 42878 60000 42880
rect 57881 42875 57947 42878
rect 59200 42788 60000 42878
rect 41597 42666 41663 42669
rect 45001 42666 45067 42669
rect 41597 42664 45067 42666
rect 41597 42608 41602 42664
rect 41658 42608 45006 42664
rect 45062 42608 45067 42664
rect 41597 42606 45067 42608
rect 41597 42603 41663 42606
rect 45001 42603 45067 42606
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 50288 42464 50608 42465
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 42399 50608 42400
rect 59200 42108 60000 42348
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 31201 41850 31267 41853
rect 34145 41850 34211 41853
rect 31201 41848 34211 41850
rect 31201 41792 31206 41848
rect 31262 41792 34150 41848
rect 34206 41792 34211 41848
rect 31201 41790 34211 41792
rect 31201 41787 31267 41790
rect 34145 41787 34211 41790
rect 20437 41714 20503 41717
rect 22553 41714 22619 41717
rect 20437 41712 22619 41714
rect 0 41428 800 41668
rect 20437 41656 20442 41712
rect 20498 41656 22558 41712
rect 22614 41656 22619 41712
rect 20437 41654 22619 41656
rect 20437 41651 20503 41654
rect 22553 41651 22619 41654
rect 20805 41578 20871 41581
rect 21909 41578 21975 41581
rect 20805 41576 21975 41578
rect 20805 41520 20810 41576
rect 20866 41520 21914 41576
rect 21970 41520 21975 41576
rect 20805 41518 21975 41520
rect 20805 41515 20871 41518
rect 21909 41515 21975 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 50288 41376 50608 41377
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 41311 50608 41312
rect 0 40748 800 40988
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 59200 40748 60000 40988
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 50288 40288 50608 40289
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 40223 50608 40224
rect 48313 39946 48379 39949
rect 53925 39946 53991 39949
rect 48313 39944 53991 39946
rect 48313 39888 48318 39944
rect 48374 39888 53930 39944
rect 53986 39888 53991 39944
rect 48313 39886 53991 39888
rect 48313 39883 48379 39886
rect 53925 39883 53991 39886
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 2773 39538 2839 39541
rect 0 39536 2839 39538
rect 0 39480 2778 39536
rect 2834 39480 2839 39536
rect 0 39478 2839 39480
rect 0 39388 800 39478
rect 2773 39475 2839 39478
rect 57881 39538 57947 39541
rect 59200 39538 60000 39628
rect 57881 39536 60000 39538
rect 57881 39480 57886 39536
rect 57942 39480 60000 39536
rect 57881 39478 60000 39480
rect 57881 39475 57947 39478
rect 59200 39388 60000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 39389 38994 39455 38997
rect 41321 38994 41387 38997
rect 39389 38992 41387 38994
rect 39389 38936 39394 38992
rect 39450 38936 41326 38992
rect 41382 38936 41387 38992
rect 39389 38934 41387 38936
rect 39389 38931 39455 38934
rect 41321 38931 41387 38934
rect 33409 38858 33475 38861
rect 34237 38858 34303 38861
rect 37089 38858 37155 38861
rect 33409 38856 37155 38858
rect 33409 38800 33414 38856
rect 33470 38800 34242 38856
rect 34298 38800 37094 38856
rect 37150 38800 37155 38856
rect 33409 38798 37155 38800
rect 33409 38795 33475 38798
rect 34237 38795 34303 38798
rect 37089 38795 37155 38798
rect 39389 38858 39455 38861
rect 40585 38858 40651 38861
rect 39389 38856 40651 38858
rect 39389 38800 39394 38856
rect 39450 38800 40590 38856
rect 40646 38800 40651 38856
rect 39389 38798 40651 38800
rect 39389 38795 39455 38798
rect 40585 38795 40651 38798
rect 57881 38858 57947 38861
rect 59200 38858 60000 38948
rect 57881 38856 60000 38858
rect 57881 38800 57886 38856
rect 57942 38800 60000 38856
rect 57881 38798 60000 38800
rect 57881 38795 57947 38798
rect 31109 38722 31175 38725
rect 31293 38722 31359 38725
rect 33593 38722 33659 38725
rect 31109 38720 33659 38722
rect 31109 38664 31114 38720
rect 31170 38664 31298 38720
rect 31354 38664 33598 38720
rect 33654 38664 33659 38720
rect 31109 38662 33659 38664
rect 31109 38659 31175 38662
rect 31293 38659 31359 38662
rect 33593 38659 33659 38662
rect 34605 38724 34671 38725
rect 34605 38720 34652 38724
rect 34716 38722 34722 38724
rect 34605 38664 34610 38720
rect 34605 38660 34652 38664
rect 34716 38662 34762 38722
rect 59200 38708 60000 38798
rect 35341 38670 35407 38673
rect 35341 38668 35450 38670
rect 34716 38660 34722 38662
rect 34605 38659 34671 38660
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 35341 38612 35346 38668
rect 35402 38612 35450 38668
rect 35341 38607 35450 38612
rect 34928 38591 35248 38592
rect 35390 38586 35450 38607
rect 41781 38586 41847 38589
rect 46381 38586 46447 38589
rect 35390 38526 35818 38586
rect 34513 38450 34579 38453
rect 35157 38450 35223 38453
rect 34513 38448 35223 38450
rect 34513 38392 34518 38448
rect 34574 38392 35162 38448
rect 35218 38392 35223 38448
rect 34513 38390 35223 38392
rect 34513 38387 34579 38390
rect 35157 38387 35223 38390
rect 30925 38314 30991 38317
rect 31293 38314 31359 38317
rect 30925 38312 31359 38314
rect 0 38028 800 38268
rect 30925 38256 30930 38312
rect 30986 38256 31298 38312
rect 31354 38256 31359 38312
rect 30925 38254 31359 38256
rect 30925 38251 30991 38254
rect 31293 38251 31359 38254
rect 34329 38314 34395 38317
rect 34513 38314 34579 38317
rect 34329 38312 34579 38314
rect 34329 38256 34334 38312
rect 34390 38256 34518 38312
rect 34574 38256 34579 38312
rect 34329 38254 34579 38256
rect 34329 38251 34395 38254
rect 34513 38251 34579 38254
rect 35341 38314 35407 38317
rect 35758 38314 35818 38526
rect 41781 38584 46447 38586
rect 41781 38528 41786 38584
rect 41842 38528 46386 38584
rect 46442 38528 46447 38584
rect 41781 38526 46447 38528
rect 41781 38523 41847 38526
rect 46381 38523 46447 38526
rect 35341 38312 35818 38314
rect 35341 38256 35346 38312
rect 35402 38256 35818 38312
rect 35341 38254 35818 38256
rect 35341 38251 35407 38254
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 39573 38042 39639 38045
rect 45277 38042 45343 38045
rect 39573 38040 45343 38042
rect 39573 37984 39578 38040
rect 39634 37984 45282 38040
rect 45338 37984 45343 38040
rect 39573 37982 45343 37984
rect 39573 37979 39639 37982
rect 45277 37979 45343 37982
rect 49785 38042 49851 38045
rect 49918 38042 49924 38044
rect 49785 38040 49924 38042
rect 49785 37984 49790 38040
rect 49846 37984 49924 38040
rect 49785 37982 49924 37984
rect 49785 37979 49851 37982
rect 49918 37980 49924 37982
rect 49988 37980 49994 38044
rect 42793 37906 42859 37909
rect 47669 37906 47735 37909
rect 42793 37904 47735 37906
rect 42793 37848 42798 37904
rect 42854 37848 47674 37904
rect 47730 37848 47735 37904
rect 42793 37846 47735 37848
rect 42793 37843 42859 37846
rect 47669 37843 47735 37846
rect 38377 37770 38443 37773
rect 40677 37770 40743 37773
rect 38377 37768 40743 37770
rect 38377 37712 38382 37768
rect 38438 37712 40682 37768
rect 40738 37712 40743 37768
rect 38377 37710 40743 37712
rect 38377 37707 38443 37710
rect 40677 37707 40743 37710
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 59200 37348 60000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 0 36668 800 36908
rect 31017 36818 31083 36821
rect 36537 36818 36603 36821
rect 37365 36818 37431 36821
rect 31017 36816 37431 36818
rect 31017 36760 31022 36816
rect 31078 36760 36542 36816
rect 36598 36760 37370 36816
rect 37426 36760 37431 36816
rect 31017 36758 37431 36760
rect 31017 36755 31083 36758
rect 36537 36755 36603 36758
rect 37365 36755 37431 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 59200 35988 60000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 42517 35186 42583 35189
rect 44265 35186 44331 35189
rect 42517 35184 44331 35186
rect 42517 35128 42522 35184
rect 42578 35128 44270 35184
rect 44326 35128 44331 35184
rect 42517 35126 44331 35128
rect 42517 35123 42583 35126
rect 44265 35123 44331 35126
rect 49877 35050 49943 35053
rect 51717 35050 51783 35053
rect 49877 35048 51783 35050
rect 49877 34992 49882 35048
rect 49938 34992 51722 35048
rect 51778 34992 51783 35048
rect 49877 34990 51783 34992
rect 49877 34987 49943 34990
rect 51717 34987 51783 34990
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 57881 34778 57947 34781
rect 59200 34778 60000 34868
rect 57881 34776 60000 34778
rect 57881 34720 57886 34776
rect 57942 34720 60000 34776
rect 57881 34718 60000 34720
rect 57881 34715 57947 34718
rect 42793 34642 42859 34645
rect 44173 34642 44239 34645
rect 42793 34640 44239 34642
rect 42793 34584 42798 34640
rect 42854 34584 44178 34640
rect 44234 34584 44239 34640
rect 42793 34582 44239 34584
rect 42793 34579 42859 34582
rect 44173 34579 44239 34582
rect 50245 34642 50311 34645
rect 51441 34642 51507 34645
rect 50245 34640 51507 34642
rect 50245 34584 50250 34640
rect 50306 34584 51446 34640
rect 51502 34584 51507 34640
rect 59200 34628 60000 34718
rect 50245 34582 51507 34584
rect 50245 34579 50311 34582
rect 51441 34579 51507 34582
rect 40401 34506 40467 34509
rect 40677 34506 40743 34509
rect 45737 34506 45803 34509
rect 40401 34504 45803 34506
rect 40401 34448 40406 34504
rect 40462 34448 40682 34504
rect 40738 34448 45742 34504
rect 45798 34448 45803 34504
rect 40401 34446 45803 34448
rect 40401 34443 40467 34446
rect 40677 34443 40743 34446
rect 45737 34443 45803 34446
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 57789 34098 57855 34101
rect 59200 34098 60000 34188
rect 57789 34096 60000 34098
rect 57789 34040 57794 34096
rect 57850 34040 60000 34096
rect 57789 34038 60000 34040
rect 57789 34035 57855 34038
rect 36077 33962 36143 33965
rect 49049 33962 49115 33965
rect 49969 33962 50035 33965
rect 36077 33960 50035 33962
rect 36077 33904 36082 33960
rect 36138 33904 49054 33960
rect 49110 33904 49974 33960
rect 50030 33904 50035 33960
rect 59200 33948 60000 34038
rect 36077 33902 50035 33904
rect 36077 33899 36143 33902
rect 49049 33899 49115 33902
rect 49969 33899 50035 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 37181 33554 37247 33557
rect 37181 33552 41430 33554
rect 0 33268 800 33508
rect 37181 33496 37186 33552
rect 37242 33496 41430 33552
rect 37181 33494 41430 33496
rect 37181 33491 37247 33494
rect 41370 33418 41430 33494
rect 49233 33418 49299 33421
rect 41370 33416 49299 33418
rect 41370 33360 49238 33416
rect 49294 33360 49299 33416
rect 41370 33358 49299 33360
rect 49233 33355 49299 33358
rect 43897 33282 43963 33285
rect 49049 33282 49115 33285
rect 43897 33280 49115 33282
rect 43897 33224 43902 33280
rect 43958 33224 49054 33280
rect 49110 33224 49115 33280
rect 43897 33222 49115 33224
rect 43897 33219 43963 33222
rect 49049 33219 49115 33222
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32588 800 32828
rect 57789 32738 57855 32741
rect 59200 32738 60000 32828
rect 57789 32736 60000 32738
rect 57789 32680 57794 32736
rect 57850 32680 60000 32736
rect 57789 32678 60000 32680
rect 57789 32675 57855 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 59200 32588 60000 32678
rect 49969 32332 50035 32333
rect 49918 32268 49924 32332
rect 49988 32330 50035 32332
rect 49988 32328 50080 32330
rect 50030 32272 50080 32328
rect 49988 32270 50080 32272
rect 49988 32268 50035 32270
rect 49969 32267 50035 32268
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31228 800 31468
rect 57881 31378 57947 31381
rect 59200 31378 60000 31468
rect 57881 31376 60000 31378
rect 57881 31320 57886 31376
rect 57942 31320 60000 31376
rect 57881 31318 60000 31320
rect 57881 31315 57947 31318
rect 59200 31228 60000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 58157 30698 58223 30701
rect 59200 30698 60000 30788
rect 58157 30696 60000 30698
rect 58157 30640 58162 30696
rect 58218 30640 60000 30696
rect 58157 30638 60000 30640
rect 58157 30635 58223 30638
rect 59200 30548 60000 30638
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 0 30018 800 30108
rect 2773 30018 2839 30021
rect 0 30016 2839 30018
rect 0 29960 2778 30016
rect 2834 29960 2839 30016
rect 0 29958 2839 29960
rect 0 29868 800 29958
rect 2773 29955 2839 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 33685 29610 33751 29613
rect 42558 29610 42564 29612
rect 33685 29608 42564 29610
rect 33685 29552 33690 29608
rect 33746 29552 42564 29608
rect 33685 29550 42564 29552
rect 33685 29547 33751 29550
rect 42558 29548 42564 29550
rect 42628 29548 42634 29612
rect 42701 29610 42767 29613
rect 43713 29610 43779 29613
rect 42701 29608 43779 29610
rect 42701 29552 42706 29608
rect 42762 29552 43718 29608
rect 43774 29552 43779 29608
rect 42701 29550 43779 29552
rect 42701 29547 42767 29550
rect 43713 29547 43779 29550
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 59200 29188 60000 29428
rect 33501 29066 33567 29069
rect 56317 29066 56383 29069
rect 33501 29064 56383 29066
rect 33501 29008 33506 29064
rect 33562 29008 56322 29064
rect 56378 29008 56383 29064
rect 33501 29006 56383 29008
rect 33501 29003 33567 29006
rect 56317 29003 56383 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3417 28658 3483 28661
rect 0 28656 3483 28658
rect 0 28600 3422 28656
rect 3478 28600 3483 28656
rect 0 28598 3483 28600
rect 0 28508 800 28598
rect 3417 28595 3483 28598
rect 40677 28386 40743 28389
rect 48037 28386 48103 28389
rect 40677 28384 48103 28386
rect 40677 28328 40682 28384
rect 40738 28328 48042 28384
rect 48098 28328 48103 28384
rect 40677 28326 48103 28328
rect 40677 28323 40743 28326
rect 48037 28323 48103 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 34053 28250 34119 28253
rect 34646 28250 34652 28252
rect 34053 28248 34652 28250
rect 34053 28192 34058 28248
rect 34114 28192 34652 28248
rect 34053 28190 34652 28192
rect 34053 28187 34119 28190
rect 34646 28188 34652 28190
rect 34716 28188 34722 28252
rect 0 27828 800 28068
rect 55213 27978 55279 27981
rect 59200 27978 60000 28068
rect 55213 27976 60000 27978
rect 55213 27920 55218 27976
rect 55274 27920 60000 27976
rect 55213 27918 60000 27920
rect 55213 27915 55279 27918
rect 31569 27842 31635 27845
rect 32121 27842 32187 27845
rect 31569 27840 32187 27842
rect 31569 27784 31574 27840
rect 31630 27784 32126 27840
rect 32182 27784 32187 27840
rect 59200 27828 60000 27918
rect 31569 27782 32187 27784
rect 31569 27779 31635 27782
rect 32121 27779 32187 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 29545 27570 29611 27573
rect 32857 27570 32923 27573
rect 29545 27568 32923 27570
rect 29545 27512 29550 27568
rect 29606 27512 32862 27568
rect 32918 27512 32923 27568
rect 29545 27510 32923 27512
rect 29545 27507 29611 27510
rect 32857 27507 32923 27510
rect 40585 27434 40651 27437
rect 42333 27434 42399 27437
rect 40585 27432 42399 27434
rect 40585 27376 40590 27432
rect 40646 27376 42338 27432
rect 42394 27376 42399 27432
rect 40585 27374 42399 27376
rect 40585 27371 40651 27374
rect 42333 27371 42399 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 0 26618 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26468 800 26558
rect 2773 26555 2839 26558
rect 58157 26618 58223 26621
rect 59200 26618 60000 26708
rect 58157 26616 60000 26618
rect 58157 26560 58162 26616
rect 58218 26560 60000 26616
rect 58157 26558 60000 26560
rect 58157 26555 58223 26558
rect 59200 26468 60000 26558
rect 30189 26346 30255 26349
rect 30741 26346 30807 26349
rect 30189 26344 30807 26346
rect 30189 26288 30194 26344
rect 30250 26288 30746 26344
rect 30802 26288 30807 26344
rect 30189 26286 30807 26288
rect 30189 26283 30255 26286
rect 30741 26283 30807 26286
rect 30925 26346 30991 26349
rect 31845 26346 31911 26349
rect 30925 26344 31911 26346
rect 30925 26288 30930 26344
rect 30986 26288 31850 26344
rect 31906 26288 31911 26344
rect 30925 26286 31911 26288
rect 30925 26283 30991 26286
rect 31845 26283 31911 26286
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 39573 25938 39639 25941
rect 40309 25938 40375 25941
rect 39573 25936 40375 25938
rect 39573 25880 39578 25936
rect 39634 25880 40314 25936
rect 40370 25880 40375 25936
rect 39573 25878 40375 25880
rect 39573 25875 39639 25878
rect 40309 25875 40375 25878
rect 58157 25938 58223 25941
rect 59200 25938 60000 26028
rect 58157 25936 60000 25938
rect 58157 25880 58162 25936
rect 58218 25880 60000 25936
rect 58157 25878 60000 25880
rect 58157 25875 58223 25878
rect 59200 25788 60000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25108 800 25348
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 40677 24850 40743 24853
rect 46381 24850 46447 24853
rect 40677 24848 46447 24850
rect 40677 24792 40682 24848
rect 40738 24792 46386 24848
rect 46442 24792 46447 24848
rect 40677 24790 46447 24792
rect 40677 24787 40743 24790
rect 46381 24787 46447 24790
rect 43621 24714 43687 24717
rect 47945 24714 48011 24717
rect 43621 24712 48011 24714
rect 0 24578 800 24668
rect 43621 24656 43626 24712
rect 43682 24656 47950 24712
rect 48006 24656 48011 24712
rect 43621 24654 48011 24656
rect 43621 24651 43687 24654
rect 47945 24651 48011 24654
rect 2773 24578 2839 24581
rect 0 24576 2839 24578
rect 0 24520 2778 24576
rect 2834 24520 2839 24576
rect 0 24518 2839 24520
rect 0 24428 800 24518
rect 2773 24515 2839 24518
rect 58157 24578 58223 24581
rect 59200 24578 60000 24668
rect 58157 24576 60000 24578
rect 58157 24520 58162 24576
rect 58218 24520 60000 24576
rect 58157 24518 60000 24520
rect 58157 24515 58223 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 59200 24428 60000 24518
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23068 800 23308
rect 59200 23068 60000 23308
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 57881 22538 57947 22541
rect 59200 22538 60000 22628
rect 57881 22536 60000 22538
rect 57881 22480 57886 22536
rect 57942 22480 60000 22536
rect 57881 22478 60000 22480
rect 57881 22475 57947 22478
rect 59200 22388 60000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21858 800 21948
rect 2773 21858 2839 21861
rect 0 21856 2839 21858
rect 0 21800 2778 21856
rect 2834 21800 2839 21856
rect 0 21798 2839 21800
rect 0 21708 800 21798
rect 2773 21795 2839 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 57789 21178 57855 21181
rect 59200 21178 60000 21268
rect 57789 21176 60000 21178
rect 57789 21120 57794 21176
rect 57850 21120 60000 21176
rect 57789 21118 60000 21120
rect 57789 21115 57855 21118
rect 59200 21028 60000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 0 20498 800 20588
rect 2773 20498 2839 20501
rect 0 20496 2839 20498
rect 0 20440 2778 20496
rect 2834 20440 2839 20496
rect 0 20438 2839 20440
rect 0 20348 800 20438
rect 2773 20435 2839 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19668 800 19908
rect 57881 19818 57947 19821
rect 59200 19818 60000 19908
rect 57881 19816 60000 19818
rect 57881 19760 57886 19816
rect 57942 19760 60000 19816
rect 57881 19758 60000 19760
rect 57881 19755 57947 19758
rect 59200 19668 60000 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 2773 18458 2839 18461
rect 0 18456 2839 18458
rect 0 18400 2778 18456
rect 2834 18400 2839 18456
rect 0 18398 2839 18400
rect 0 18308 800 18398
rect 2773 18395 2839 18398
rect 59200 18308 60000 18548
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 58157 17778 58223 17781
rect 59200 17778 60000 17868
rect 58157 17776 60000 17778
rect 58157 17720 58162 17776
rect 58218 17720 60000 17776
rect 58157 17718 60000 17720
rect 58157 17715 58223 17718
rect 59200 17628 60000 17718
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 0 17098 800 17188
rect 2773 17098 2839 17101
rect 0 17096 2839 17098
rect 0 17040 2778 17096
rect 2834 17040 2839 17096
rect 0 17038 2839 17040
rect 0 16948 800 17038
rect 2773 17035 2839 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16268 800 16508
rect 57789 16418 57855 16421
rect 59200 16418 60000 16508
rect 57789 16416 60000 16418
rect 57789 16360 57794 16416
rect 57850 16360 60000 16416
rect 57789 16358 60000 16360
rect 57789 16355 57855 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 59200 16268 60000 16358
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 0 14908 800 15148
rect 57881 15058 57947 15061
rect 59200 15058 60000 15148
rect 57881 15056 60000 15058
rect 57881 15000 57886 15056
rect 57942 15000 60000 15056
rect 57881 14998 60000 15000
rect 57881 14995 57947 14998
rect 59200 14908 60000 14998
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 58157 14378 58223 14381
rect 59200 14378 60000 14468
rect 58157 14376 60000 14378
rect 58157 14320 58162 14376
rect 58218 14320 60000 14376
rect 58157 14318 60000 14320
rect 58157 14315 58223 14318
rect 59200 14228 60000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 0 13698 800 13788
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13548 800 13638
rect 2773 13635 2839 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 59200 12868 60000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 3969 12338 4035 12341
rect 0 12336 4035 12338
rect 0 12280 3974 12336
rect 4030 12280 4035 12336
rect 0 12278 4035 12280
rect 0 12188 800 12278
rect 3969 12275 4035 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 0 11658 800 11748
rect 2773 11658 2839 11661
rect 0 11656 2839 11658
rect 0 11600 2778 11656
rect 2834 11600 2839 11656
rect 0 11598 2839 11600
rect 0 11508 800 11598
rect 2773 11595 2839 11598
rect 59200 11508 60000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 0 10148 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 59200 10148 60000 10388
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 57237 9618 57303 9621
rect 59200 9618 60000 9708
rect 57237 9616 60000 9618
rect 57237 9560 57242 9616
rect 57298 9560 60000 9616
rect 57237 9558 60000 9560
rect 57237 9555 57303 9558
rect 59200 9468 60000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 9028
rect 3417 8938 3483 8941
rect 0 8936 3483 8938
rect 0 8880 3422 8936
rect 3478 8880 3483 8936
rect 0 8878 3483 8880
rect 0 8788 800 8878
rect 3417 8875 3483 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 0 8258 800 8348
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8108 800 8198
rect 2773 8195 2839 8198
rect 57881 8258 57947 8261
rect 59200 8258 60000 8348
rect 57881 8256 60000 8258
rect 57881 8200 57886 8256
rect 57942 8200 60000 8256
rect 57881 8198 60000 8200
rect 57881 8195 57947 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 59200 8108 60000 8198
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6748 800 6838
rect 2773 6835 2839 6838
rect 59200 6748 60000 6988
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 58157 6218 58223 6221
rect 59200 6218 60000 6308
rect 58157 6216 60000 6218
rect 58157 6160 58162 6216
rect 58218 6160 60000 6216
rect 58157 6158 60000 6160
rect 58157 6155 58223 6158
rect 59200 6068 60000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5538 800 5628
rect 3233 5538 3299 5541
rect 0 5536 3299 5538
rect 0 5480 3238 5536
rect 3294 5480 3299 5536
rect 0 5478 3299 5480
rect 0 5388 800 5478
rect 3233 5475 3299 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 59200 4708 60000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 0 4178 800 4268
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4028 800 4118
rect 2773 4115 2839 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 2865 3498 2931 3501
rect 0 3496 2931 3498
rect 0 3440 2870 3496
rect 2926 3440 2931 3496
rect 0 3438 2931 3440
rect 0 3348 800 3438
rect 2865 3435 2931 3438
rect 59200 3348 60000 3588
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 0 2138 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 1988 800 2078
rect 2773 2075 2839 2078
rect 57697 2138 57763 2141
rect 59200 2138 60000 2228
rect 57697 2136 60000 2138
rect 57697 2080 57702 2136
rect 57758 2080 60000 2136
rect 57697 2078 60000 2080
rect 57697 2075 57763 2078
rect 59200 1988 60000 2078
rect 57881 1458 57947 1461
rect 59200 1458 60000 1548
rect 57881 1456 60000 1458
rect 57881 1400 57886 1456
rect 57942 1400 60000 1456
rect 57881 1398 60000 1400
rect 57881 1395 57947 1398
rect 59200 1308 60000 1398
rect 0 628 800 868
rect 56501 98 56567 101
rect 59200 98 60000 188
rect 56501 96 60000 98
rect 56501 40 56506 96
rect 56562 40 60000 96
rect 56501 38 60000 40
rect 56501 35 56567 38
rect 59200 -52 60000 38
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 42564 55448 42628 55452
rect 42564 55392 42614 55448
rect 42614 55392 42628 55448
rect 42564 55388 42628 55392
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 34652 38720 34716 38724
rect 34652 38664 34666 38720
rect 34666 38664 34716 38720
rect 34652 38660 34716 38664
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 49924 37980 49988 38044
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 49924 32328 49988 32332
rect 49924 32272 49974 32328
rect 49974 32272 49988 32328
rect 49924 32268 49988 32272
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 42564 29548 42628 29612
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 34652 28188 34716 28252
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 42563 55452 42629 55453
rect 42563 55388 42564 55452
rect 42628 55388 42629 55452
rect 42563 55387 42629 55388
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34651 38724 34717 38725
rect 34651 38660 34652 38724
rect 34716 38660 34717 38724
rect 34651 38659 34717 38660
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 34654 28253 34714 38659
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 42566 29613 42626 55387
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 49923 38044 49989 38045
rect 49923 37980 49924 38044
rect 49988 37980 49989 38044
rect 49923 37979 49989 37980
rect 49926 32333 49986 37979
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 49923 32332 49989 32333
rect 49923 32268 49924 32332
rect 49988 32268 49989 32332
rect 49923 32267 49989 32268
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 42563 29612 42629 29613
rect 42563 29548 42564 29612
rect 42628 29548 42629 29612
rect 42563 29547 42629 29548
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34651 28252 34717 28253
rect 34651 28188 34652 28252
rect 34716 28188 34717 28252
rect 34651 28187 34717 28188
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 20424 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_325
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1644511149
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1644511149
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1644511149
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_517
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_561
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1644511149
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1644511149
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1644511149
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1644511149
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1644511149
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_36
timestamp 1644511149
transform 1 0 4416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_64
timestamp 1644511149
transform 1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_145
timestamp 1644511149
transform 1 0 14444 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_156
timestamp 1644511149
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_202
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_212
timestamp 1644511149
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1644511149
transform 1 0 24748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1644511149
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_296
timestamp 1644511149
transform 1 0 28336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_308
timestamp 1644511149
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_341
timestamp 1644511149
transform 1 0 32476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_357
timestamp 1644511149
transform 1 0 33948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_369
timestamp 1644511149
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_381
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp 1644511149
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_401
timestamp 1644511149
transform 1 0 37996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_425
timestamp 1644511149
transform 1 0 40204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_437
timestamp 1644511149
transform 1 0 41308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_445
timestamp 1644511149
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_493
timestamp 1644511149
transform 1 0 46460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_499
timestamp 1644511149
transform 1 0 47012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_533
timestamp 1644511149
transform 1 0 50140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_545
timestamp 1644511149
transform 1 0 51244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1644511149
transform 1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_567
timestamp 1644511149
transform 1 0 53268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1644511149
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_596
timestamp 1644511149
transform 1 0 55936 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_604
timestamp 1644511149
transform 1 0 56672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1644511149
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1644511149
transform 1 0 58512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1644511149
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1644511149
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_111
timestamp 1644511149
transform 1 0 11316 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_119
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1644511149
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_131
timestamp 1644511149
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_149
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1644511149
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_205
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_230
timestamp 1644511149
transform 1 0 22264 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_239
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_274
timestamp 1644511149
transform 1 0 26312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 1644511149
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1644511149
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_408
timestamp 1644511149
transform 1 0 38640 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_519
timestamp 1644511149
transform 1 0 48852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_528
timestamp 1644511149
transform 1 0 49680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_554
timestamp 1644511149
transform 1 0 52072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_562
timestamp 1644511149
transform 1 0 52808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1644511149
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_592
timestamp 1644511149
transform 1 0 55568 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_40
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_96
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1644511149
transform 1 0 19136 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp 1644511149
transform 1 0 22356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_254
timestamp 1644511149
transform 1 0 24472 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_266
timestamp 1644511149
transform 1 0 25576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1644511149
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_284
timestamp 1644511149
transform 1 0 27232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_296
timestamp 1644511149
transform 1 0 28336 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_308
timestamp 1644511149
transform 1 0 29440 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_315
timestamp 1644511149
transform 1 0 30084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_322
timestamp 1644511149
transform 1 0 30728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_340
timestamp 1644511149
transform 1 0 32384 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_352
timestamp 1644511149
transform 1 0 33488 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_364
timestamp 1644511149
transform 1 0 34592 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_376
timestamp 1644511149
transform 1 0 35696 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_404
timestamp 1644511149
transform 1 0 38272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_416
timestamp 1644511149
transform 1 0 39376 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_428
timestamp 1644511149
transform 1 0 40480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1644511149
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_494
timestamp 1644511149
transform 1 0 46552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1644511149
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_534
timestamp 1644511149
transform 1 0 50232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_546
timestamp 1644511149
transform 1 0 51336 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_558
timestamp 1644511149
transform 1 0 52440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_576
timestamp 1644511149
transform 1 0 54096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_587
timestamp 1644511149
transform 1 0 55108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_612
timestamp 1644511149
transform 1 0 57408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_620
timestamp 1644511149
transform 1 0 58144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_624
timestamp 1644511149
transform 1 0 58512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1644511149
transform 1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_16
timestamp 1644511149
transform 1 0 2576 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_90
timestamp 1644511149
transform 1 0 9384 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_102
timestamp 1644511149
transform 1 0 10488 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_114
timestamp 1644511149
transform 1 0 11592 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_126
timestamp 1644511149
transform 1 0 12696 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1644511149
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_584
timestamp 1644511149
transform 1 0 54832 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_596
timestamp 1644511149
transform 1 0 55936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1644511149
transform 1 0 58236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1644511149
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp 1644511149
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_79
timestamp 1644511149
transform 1 0 8372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_91
timestamp 1644511149
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_612
timestamp 1644511149
transform 1 0 57408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_620
timestamp 1644511149
transform 1 0 58144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_624
timestamp 1644511149
transform 1 0 58512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1644511149
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_16
timestamp 1644511149
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_596
timestamp 1644511149
transform 1 0 55936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1644511149
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1644511149
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_591
timestamp 1644511149
transform 1 0 55476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_612
timestamp 1644511149
transform 1 0 57408 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_620
timestamp 1644511149
transform 1 0 58144 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_624
timestamp 1644511149
transform 1 0 58512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1644511149
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1644511149
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1644511149
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1644511149
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_610
timestamp 1644511149
transform 1 0 57224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_617
timestamp 1644511149
transform 1 0 57868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1644511149
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_37
timestamp 1644511149
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1644511149
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1644511149
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1644511149
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1644511149
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1644511149
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_597
timestamp 1644511149
transform 1 0 56028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1644511149
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_312
timestamp 1644511149
transform 1 0 29808 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_324
timestamp 1644511149
transform 1 0 30912 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_620
timestamp 1644511149
transform 1 0 58144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_624
timestamp 1644511149
transform 1 0 58512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_330
timestamp 1644511149
transform 1 0 31464 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_342
timestamp 1644511149
transform 1 0 32568 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_354
timestamp 1644511149
transform 1 0 33672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1644511149
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_606
timestamp 1644511149
transform 1 0 56856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1644511149
transform 1 0 58236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_16
timestamp 1644511149
transform 1 0 2576 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_30
timestamp 1644511149
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_42
timestamp 1644511149
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1644511149
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1644511149
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_13
timestamp 1644511149
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1644511149
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1644511149
transform 1 0 4048 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1644511149
transform 1 0 5152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1644511149
transform 1 0 6256 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1644511149
transform 1 0 7360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_8
timestamp 1644511149
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_33
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1644511149
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_11
timestamp 1644511149
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_17
timestamp 1644511149
transform 1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1644511149
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_30
timestamp 1644511149
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_42
timestamp 1644511149
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1644511149
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_605
timestamp 1644511149
transform 1 0 56764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1644511149
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_13
timestamp 1644511149
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1644511149
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_597
timestamp 1644511149
transform 1 0 56028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1644511149
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_605
timestamp 1644511149
transform 1 0 56764 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_620
timestamp 1644511149
transform 1 0 58144 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_624
timestamp 1644511149
transform 1 0 58512 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_597
timestamp 1644511149
transform 1 0 56028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_621
timestamp 1644511149
transform 1 0 58236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_605
timestamp 1644511149
transform 1 0 56764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_611
timestamp 1644511149
transform 1 0 57316 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_620
timestamp 1644511149
transform 1 0 58144 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_624
timestamp 1644511149
transform 1 0 58512 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_16
timestamp 1644511149
transform 1 0 2576 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_597
timestamp 1644511149
transform 1 0 56028 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1644511149
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_30
timestamp 1644511149
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_42
timestamp 1644511149
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1644511149
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_605
timestamp 1644511149
transform 1 0 56764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_611
timestamp 1644511149
transform 1 0 57316 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_620
timestamp 1644511149
transform 1 0 58144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_624
timestamp 1644511149
transform 1 0 58512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1644511149
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_13
timestamp 1644511149
transform 1 0 2300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1644511149
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_346
timestamp 1644511149
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1644511149
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_597
timestamp 1644511149
transform 1 0 56028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_621
timestamp 1644511149
transform 1 0 58236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_33
timestamp 1644511149
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1644511149
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1644511149
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_321
timestamp 1644511149
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1644511149
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_620
timestamp 1644511149
transform 1 0 58144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_624
timestamp 1644511149
transform 1 0 58512 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_16
timestamp 1644511149
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1644511149
transform 1 0 4048 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1644511149
transform 1 0 5152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1644511149
transform 1 0 6256 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1644511149
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1644511149
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1644511149
transform 1 0 2668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1644511149
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1644511149
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1644511149
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_315
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_327
timestamp 1644511149
transform 1 0 31188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1644511149
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1644511149
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_216
timestamp 1644511149
transform 1 0 20976 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_228
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_240
timestamp 1644511149
transform 1 0 23184 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_317
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_331
timestamp 1644511149
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_343
timestamp 1644511149
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1644511149
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_597
timestamp 1644511149
transform 1 0 56028 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1644511149
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_30
timestamp 1644511149
transform 1 0 3864 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_42
timestamp 1644511149
transform 1 0 4968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1644511149
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1644511149
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_309
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_326
timestamp 1644511149
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1644511149
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_620
timestamp 1644511149
transform 1 0 58144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_624
timestamp 1644511149
transform 1 0 58512 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1644511149
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_13
timestamp 1644511149
transform 1 0 2300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1644511149
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_185
timestamp 1644511149
transform 1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_297
timestamp 1644511149
transform 1 0 28428 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_317
timestamp 1644511149
transform 1 0 30268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_331
timestamp 1644511149
transform 1 0 31556 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_343
timestamp 1644511149
transform 1 0 32660 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_355
timestamp 1644511149
transform 1 0 33764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_597
timestamp 1644511149
transform 1 0 56028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_621
timestamp 1644511149
transform 1 0 58236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_30
timestamp 1644511149
transform 1 0 3864 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1644511149
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1644511149
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_176
timestamp 1644511149
transform 1 0 17296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_188
timestamp 1644511149
transform 1 0 18400 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_209
timestamp 1644511149
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1644511149
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 1644511149
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_605
timestamp 1644511149
transform 1 0 56764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_610
timestamp 1644511149
transform 1 0 57224 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_620
timestamp 1644511149
transform 1 0 58144 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_624
timestamp 1644511149
transform 1 0 58512 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1644511149
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_13
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_25
timestamp 1644511149
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_464
timestamp 1644511149
transform 1 0 43792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1644511149
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_597
timestamp 1644511149
transform 1 0 56028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_621
timestamp 1644511149
transform 1 0 58236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_457
timestamp 1644511149
transform 1 0 43148 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_464
timestamp 1644511149
transform 1 0 43792 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_475
timestamp 1644511149
transform 1 0 44804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_482
timestamp 1644511149
transform 1 0 45448 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_494
timestamp 1644511149
transform 1 0 46552 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1644511149
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_601
timestamp 1644511149
transform 1 0 56396 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_605
timestamp 1644511149
transform 1 0 56764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_612
timestamp 1644511149
transform 1 0 57408 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_620
timestamp 1644511149
transform 1 0 58144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_624
timestamp 1644511149
transform 1 0 58512 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_428
timestamp 1644511149
transform 1 0 40480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_439
timestamp 1644511149
transform 1 0 41492 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_449
timestamp 1644511149
transform 1 0 42412 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_465
timestamp 1644511149
transform 1 0 43884 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1644511149
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_486
timestamp 1644511149
transform 1 0 45816 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_30
timestamp 1644511149
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_42
timestamp 1644511149
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1644511149
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_344
timestamp 1644511149
transform 1 0 32752 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_356
timestamp 1644511149
transform 1 0 33856 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_368
timestamp 1644511149
transform 1 0 34960 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_380
timestamp 1644511149
transform 1 0 36064 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_457
timestamp 1644511149
transform 1 0 43148 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_463
timestamp 1644511149
transform 1 0 43700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_475
timestamp 1644511149
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_486
timestamp 1644511149
transform 1 0 45816 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_499
timestamp 1644511149
transform 1 0 47012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_510
timestamp 1644511149
transform 1 0 48024 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_522
timestamp 1644511149
transform 1 0 49128 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_534
timestamp 1644511149
transform 1 0 50232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_546
timestamp 1644511149
transform 1 0 51336 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_558
timestamp 1644511149
transform 1 0 52440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_427
timestamp 1644511149
transform 1 0 40388 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_435
timestamp 1644511149
transform 1 0 41124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_444
timestamp 1644511149
transform 1 0 41952 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_450
timestamp 1644511149
transform 1 0 42504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_456
timestamp 1644511149
transform 1 0 43056 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_464
timestamp 1644511149
transform 1 0 43792 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_472
timestamp 1644511149
transform 1 0 44528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_485
timestamp 1644511149
transform 1 0 45724 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_504
timestamp 1644511149
transform 1 0 47472 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_515
timestamp 1644511149
transform 1 0 48484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_523
timestamp 1644511149
transform 1 0 49220 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_597
timestamp 1644511149
transform 1 0 56028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1644511149
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1644511149
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_16
timestamp 1644511149
transform 1 0 2576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_28
timestamp 1644511149
transform 1 0 3680 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_40
timestamp 1644511149
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1644511149
transform 1 0 9752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1644511149
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_398
timestamp 1644511149
transform 1 0 37720 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_410
timestamp 1644511149
transform 1 0 38824 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_419
timestamp 1644511149
transform 1 0 39652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_430
timestamp 1644511149
transform 1 0 40664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_455
timestamp 1644511149
transform 1 0 42964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_463
timestamp 1644511149
transform 1 0 43700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_476
timestamp 1644511149
transform 1 0 44896 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_486
timestamp 1644511149
transform 1 0 45816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_490
timestamp 1644511149
transform 1 0 46184 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_511
timestamp 1644511149
transform 1 0 48116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_523
timestamp 1644511149
transform 1 0 49220 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_535
timestamp 1644511149
transform 1 0 50324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_547
timestamp 1644511149
transform 1 0 51428 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_605
timestamp 1644511149
transform 1 0 56764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_620
timestamp 1644511149
transform 1 0 58144 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_624
timestamp 1644511149
transform 1 0 58512 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_113
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1644511149
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_381
timestamp 1644511149
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_400
timestamp 1644511149
transform 1 0 37904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_407
timestamp 1644511149
transform 1 0 38548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1644511149
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_428
timestamp 1644511149
transform 1 0 40480 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_436
timestamp 1644511149
transform 1 0 41216 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_440
timestamp 1644511149
transform 1 0 41584 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_465
timestamp 1644511149
transform 1 0 43884 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_472
timestamp 1644511149
transform 1 0 44528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_481
timestamp 1644511149
transform 1 0 45356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_493
timestamp 1644511149
transform 1 0 46460 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_499
timestamp 1644511149
transform 1 0 47012 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_503
timestamp 1644511149
transform 1 0 47380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_510
timestamp 1644511149
transform 1 0 48024 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_522
timestamp 1644511149
transform 1 0 49128 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_530
timestamp 1644511149
transform 1 0 49864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_597
timestamp 1644511149
transform 1 0 56028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1644511149
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_77
timestamp 1644511149
transform 1 0 8188 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_97
timestamp 1644511149
transform 1 0 10028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1644511149
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_313
timestamp 1644511149
transform 1 0 29900 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_323
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_330
timestamp 1644511149
transform 1 0 31464 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_414
timestamp 1644511149
transform 1 0 39192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_426
timestamp 1644511149
transform 1 0 40296 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_434
timestamp 1644511149
transform 1 0 41032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_444
timestamp 1644511149
transform 1 0 41952 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_457
timestamp 1644511149
transform 1 0 43148 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_465
timestamp 1644511149
transform 1 0 43884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_476
timestamp 1644511149
transform 1 0 44896 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_488
timestamp 1644511149
transform 1 0 46000 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1644511149
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_524
timestamp 1644511149
transform 1 0 49312 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_536
timestamp 1644511149
transform 1 0 50416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_548
timestamp 1644511149
transform 1 0 51520 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_603
timestamp 1644511149
transform 1 0 56580 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_610
timestamp 1644511149
transform 1 0 57224 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_620
timestamp 1644511149
transform 1 0 58144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_624
timestamp 1644511149
transform 1 0 58512 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_17
timestamp 1644511149
transform 1 0 2668 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1644511149
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_314
timestamp 1644511149
transform 1 0 29992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_327
timestamp 1644511149
transform 1 0 31188 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_338
timestamp 1644511149
transform 1 0 32200 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_350
timestamp 1644511149
transform 1 0 33304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1644511149
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_393
timestamp 1644511149
transform 1 0 37260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_400
timestamp 1644511149
transform 1 0 37904 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_412
timestamp 1644511149
transform 1 0 39008 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_427
timestamp 1644511149
transform 1 0 40388 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_434
timestamp 1644511149
transform 1 0 41032 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_441
timestamp 1644511149
transform 1 0 41676 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_453
timestamp 1644511149
transform 1 0 42780 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_460
timestamp 1644511149
transform 1 0 43424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_472
timestamp 1644511149
transform 1 0 44528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_497
timestamp 1644511149
transform 1 0 46828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_504
timestamp 1644511149
transform 1 0 47472 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_511
timestamp 1644511149
transform 1 0 48116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_523
timestamp 1644511149
transform 1 0 49220 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_539
timestamp 1644511149
transform 1 0 50692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_548
timestamp 1644511149
transform 1 0 51520 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_560
timestamp 1644511149
transform 1 0 52624 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_572
timestamp 1644511149
transform 1 0 53728 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_584
timestamp 1644511149
transform 1 0 54832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_597
timestamp 1644511149
transform 1 0 56028 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_621
timestamp 1644511149
transform 1 0 58236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_30
timestamp 1644511149
transform 1 0 3864 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_42
timestamp 1644511149
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1644511149
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_91
timestamp 1644511149
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_103
timestamp 1644511149
transform 1 0 10580 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_302
timestamp 1644511149
transform 1 0 28888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_309
timestamp 1644511149
transform 1 0 29532 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_323
timestamp 1644511149
transform 1 0 30820 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_343
timestamp 1644511149
transform 1 0 32660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_355
timestamp 1644511149
transform 1 0 33764 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1644511149
transform 1 0 34868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_379
timestamp 1644511149
transform 1 0 35972 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1644511149
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_400
timestamp 1644511149
transform 1 0 37904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_412
timestamp 1644511149
transform 1 0 39008 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_420
timestamp 1644511149
transform 1 0 39744 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_427
timestamp 1644511149
transform 1 0 40388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_431
timestamp 1644511149
transform 1 0 40756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_442
timestamp 1644511149
transform 1 0 41768 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_466
timestamp 1644511149
transform 1 0 43976 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_478
timestamp 1644511149
transform 1 0 45080 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_490
timestamp 1644511149
transform 1 0 46184 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_500
timestamp 1644511149
transform 1 0 47104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_515
timestamp 1644511149
transform 1 0 48484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_524
timestamp 1644511149
transform 1 0 49312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_538
timestamp 1644511149
transform 1 0 50600 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_552
timestamp 1644511149
transform 1 0 51888 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_605
timestamp 1644511149
transform 1 0 56764 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_610
timestamp 1644511149
transform 1 0 57224 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_620
timestamp 1644511149
transform 1 0 58144 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_624
timestamp 1644511149
transform 1 0 58512 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1644511149
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1644511149
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_326
timestamp 1644511149
transform 1 0 31096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_337
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_346
timestamp 1644511149
transform 1 0 32936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_353
timestamp 1644511149
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1644511149
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_384
timestamp 1644511149
transform 1 0 36432 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_394
timestamp 1644511149
transform 1 0 37352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1644511149
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_411
timestamp 1644511149
transform 1 0 38916 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_431
timestamp 1644511149
transform 1 0 40756 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_443
timestamp 1644511149
transform 1 0 41860 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_451
timestamp 1644511149
transform 1 0 42596 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_459
timestamp 1644511149
transform 1 0 43332 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_467
timestamp 1644511149
transform 1 0 44068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_483
timestamp 1644511149
transform 1 0 45540 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_493
timestamp 1644511149
transform 1 0 46460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_505
timestamp 1644511149
transform 1 0 47564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_516
timestamp 1644511149
transform 1 0 48576 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_520
timestamp 1644511149
transform 1 0 48944 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_528
timestamp 1644511149
transform 1 0 49680 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_543
timestamp 1644511149
transform 1 0 51060 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_565
timestamp 1644511149
transform 1 0 53084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_572
timestamp 1644511149
transform 1 0 53728 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_584
timestamp 1644511149
transform 1 0 54832 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_605
timestamp 1644511149
transform 1 0 56764 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_609
timestamp 1644511149
transform 1 0 57132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_621
timestamp 1644511149
transform 1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_301
timestamp 1644511149
transform 1 0 28796 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_306
timestamp 1644511149
transform 1 0 29256 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_316
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_343
timestamp 1644511149
transform 1 0 32660 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_351
timestamp 1644511149
transform 1 0 33396 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_372
timestamp 1644511149
transform 1 0 35328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_379
timestamp 1644511149
transform 1 0 35972 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_410
timestamp 1644511149
transform 1 0 38824 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_437
timestamp 1644511149
transform 1 0 41308 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_445
timestamp 1644511149
transform 1 0 42044 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_460
timestamp 1644511149
transform 1 0 43424 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_471
timestamp 1644511149
transform 1 0 44436 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_478
timestamp 1644511149
transform 1 0 45080 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_489
timestamp 1644511149
transform 1 0 46092 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_496
timestamp 1644511149
transform 1 0 46736 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_510
timestamp 1644511149
transform 1 0 48024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_522
timestamp 1644511149
transform 1 0 49128 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_528
timestamp 1644511149
transform 1 0 49680 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_542
timestamp 1644511149
transform 1 0 50968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_569
timestamp 1644511149
transform 1 0 53452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_576
timestamp 1644511149
transform 1 0 54096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_583
timestamp 1644511149
transform 1 0 54740 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_595
timestamp 1644511149
transform 1 0 55844 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_607
timestamp 1644511149
transform 1 0 56948 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_620
timestamp 1644511149
transform 1 0 58144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_624
timestamp 1644511149
transform 1 0 58512 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_264
timestamp 1644511149
transform 1 0 25392 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_276
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_282
timestamp 1644511149
transform 1 0 27048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_286
timestamp 1644511149
transform 1 0 27416 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_319
timestamp 1644511149
transform 1 0 30452 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_327
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_338
timestamp 1644511149
transform 1 0 32200 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_347
timestamp 1644511149
transform 1 0 33028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_354
timestamp 1644511149
transform 1 0 33672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1644511149
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_382
timestamp 1644511149
transform 1 0 36248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_390
timestamp 1644511149
transform 1 0 36984 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_402
timestamp 1644511149
transform 1 0 38088 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_408
timestamp 1644511149
transform 1 0 38640 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_431
timestamp 1644511149
transform 1 0 40756 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_439
timestamp 1644511149
transform 1 0 41492 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_451
timestamp 1644511149
transform 1 0 42596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_466
timestamp 1644511149
transform 1 0 43976 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_474
timestamp 1644511149
transform 1 0 44712 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_485
timestamp 1644511149
transform 1 0 45724 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_499
timestamp 1644511149
transform 1 0 47012 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_509
timestamp 1644511149
transform 1 0 47932 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_519
timestamp 1644511149
transform 1 0 48852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_543
timestamp 1644511149
transform 1 0 51060 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_552
timestamp 1644511149
transform 1 0 51888 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_564
timestamp 1644511149
transform 1 0 52992 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_572
timestamp 1644511149
transform 1 0 53728 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_583
timestamp 1644511149
transform 1 0 54740 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_597
timestamp 1644511149
transform 1 0 56028 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_621
timestamp 1644511149
transform 1 0 58236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_30
timestamp 1644511149
transform 1 0 3864 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_42
timestamp 1644511149
transform 1 0 4968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1644511149
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_298
timestamp 1644511149
transform 1 0 28520 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_310
timestamp 1644511149
transform 1 0 29624 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_318
timestamp 1644511149
transform 1 0 30360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_327
timestamp 1644511149
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_342
timestamp 1644511149
transform 1 0 32568 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_348
timestamp 1644511149
transform 1 0 33120 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_353
timestamp 1644511149
transform 1 0 33580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_365
timestamp 1644511149
transform 1 0 34684 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_377
timestamp 1644511149
transform 1 0 35788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1644511149
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_398
timestamp 1644511149
transform 1 0 37720 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_412
timestamp 1644511149
transform 1 0 39008 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_426
timestamp 1644511149
transform 1 0 40296 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_433
timestamp 1644511149
transform 1 0 40940 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_445
timestamp 1644511149
transform 1 0 42044 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_453
timestamp 1644511149
transform 1 0 42780 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_464
timestamp 1644511149
transform 1 0 43792 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_476
timestamp 1644511149
transform 1 0 44896 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_484
timestamp 1644511149
transform 1 0 45632 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_490
timestamp 1644511149
transform 1 0 46184 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_502
timestamp 1644511149
transform 1 0 47288 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_533
timestamp 1644511149
transform 1 0 50140 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_537
timestamp 1644511149
transform 1 0 50508 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_545
timestamp 1644511149
transform 1 0 51244 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_555
timestamp 1644511149
transform 1 0 52164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_568
timestamp 1644511149
transform 1 0 53360 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_581
timestamp 1644511149
transform 1 0 54556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_593
timestamp 1644511149
transform 1 0 55660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_605
timestamp 1644511149
transform 1 0 56764 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_613
timestamp 1644511149
transform 1 0 57500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_296
timestamp 1644511149
transform 1 0 28336 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_328
timestamp 1644511149
transform 1 0 31280 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_336
timestamp 1644511149
transform 1 0 32016 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_348
timestamp 1644511149
transform 1 0 33120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_352
timestamp 1644511149
transform 1 0 33488 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1644511149
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_383
timestamp 1644511149
transform 1 0 36340 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_397
timestamp 1644511149
transform 1 0 37628 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1644511149
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_415
timestamp 1644511149
transform 1 0 39284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_428
timestamp 1644511149
transform 1 0 40480 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_436
timestamp 1644511149
transform 1 0 41216 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_442
timestamp 1644511149
transform 1 0 41768 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_450
timestamp 1644511149
transform 1 0 42504 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_458
timestamp 1644511149
transform 1 0 43240 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_468
timestamp 1644511149
transform 1 0 44160 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_480
timestamp 1644511149
transform 1 0 45264 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_499
timestamp 1644511149
transform 1 0 47012 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_510
timestamp 1644511149
transform 1 0 48024 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_522
timestamp 1644511149
transform 1 0 49128 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_530
timestamp 1644511149
transform 1 0 49864 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_548
timestamp 1644511149
transform 1 0 51520 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_556
timestamp 1644511149
transform 1 0 52256 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_567
timestamp 1644511149
transform 1 0 53268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_592
timestamp 1644511149
transform 1 0 55568 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_621
timestamp 1644511149
transform 1 0 58236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_10
timestamp 1644511149
transform 1 0 2024 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_17
timestamp 1644511149
transform 1 0 2668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_29
timestamp 1644511149
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_41
timestamp 1644511149
transform 1 0 4876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1644511149
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_269
timestamp 1644511149
transform 1 0 25852 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1644511149
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_309
timestamp 1644511149
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_327
timestamp 1644511149
transform 1 0 31188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_355
timestamp 1644511149
transform 1 0 33764 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_381
timestamp 1644511149
transform 1 0 36156 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1644511149
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_399
timestamp 1644511149
transform 1 0 37812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_411
timestamp 1644511149
transform 1 0 38916 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_418
timestamp 1644511149
transform 1 0 39560 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_437
timestamp 1644511149
transform 1 0 41308 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_444
timestamp 1644511149
transform 1 0 41952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_454
timestamp 1644511149
transform 1 0 42872 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_463
timestamp 1644511149
transform 1 0 43700 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_471
timestamp 1644511149
transform 1 0 44436 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_481
timestamp 1644511149
transform 1 0 45356 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_493
timestamp 1644511149
transform 1 0 46460 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_501
timestamp 1644511149
transform 1 0 47196 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_509
timestamp 1644511149
transform 1 0 47932 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_521
timestamp 1644511149
transform 1 0 49036 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_528
timestamp 1644511149
transform 1 0 49680 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_550
timestamp 1644511149
transform 1 0 51704 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_558
timestamp 1644511149
transform 1 0 52440 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_586
timestamp 1644511149
transform 1 0 55016 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_595
timestamp 1644511149
transform 1 0 55844 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_607
timestamp 1644511149
transform 1 0 56948 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_612
timestamp 1644511149
transform 1 0 57408 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_620
timestamp 1644511149
transform 1 0 58144 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_624
timestamp 1644511149
transform 1 0 58512 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_285
timestamp 1644511149
transform 1 0 27324 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_290
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_294
timestamp 1644511149
transform 1 0 28152 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_341
timestamp 1644511149
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_353
timestamp 1644511149
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1644511149
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_373
timestamp 1644511149
transform 1 0 35420 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_380
timestamp 1644511149
transform 1 0 36064 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_392
timestamp 1644511149
transform 1 0 37168 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_400
timestamp 1644511149
transform 1 0 37904 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_408
timestamp 1644511149
transform 1 0 38640 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1644511149
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_432
timestamp 1644511149
transform 1 0 40848 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_439
timestamp 1644511149
transform 1 0 41492 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_451
timestamp 1644511149
transform 1 0 42596 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_459
timestamp 1644511149
transform 1 0 43332 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_463
timestamp 1644511149
transform 1 0 43700 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_472
timestamp 1644511149
transform 1 0 44528 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_487
timestamp 1644511149
transform 1 0 45908 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_497
timestamp 1644511149
transform 1 0 46828 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_509
timestamp 1644511149
transform 1 0 47932 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_514
timestamp 1644511149
transform 1 0 48392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_518
timestamp 1644511149
transform 1 0 48760 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_541
timestamp 1644511149
transform 1 0 50876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_550
timestamp 1644511149
transform 1 0 51704 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_559
timestamp 1644511149
transform 1 0 52532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_571
timestamp 1644511149
transform 1 0 53636 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_579
timestamp 1644511149
transform 1 0 54372 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_583
timestamp 1644511149
transform 1 0 54740 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_595
timestamp 1644511149
transform 1 0 55844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_599
timestamp 1644511149
transform 1 0 56212 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_621
timestamp 1644511149
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_257
timestamp 1644511149
transform 1 0 24748 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_263
timestamp 1644511149
transform 1 0 25300 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1644511149
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_292
timestamp 1644511149
transform 1 0 27968 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_313
timestamp 1644511149
transform 1 0 29900 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_319
timestamp 1644511149
transform 1 0 30452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_346
timestamp 1644511149
transform 1 0 32936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_358
timestamp 1644511149
transform 1 0 34040 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_366
timestamp 1644511149
transform 1 0 34776 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_384
timestamp 1644511149
transform 1 0 36432 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_409
timestamp 1644511149
transform 1 0 38732 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_423
timestamp 1644511149
transform 1 0 40020 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_430
timestamp 1644511149
transform 1 0 40664 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_442
timestamp 1644511149
transform 1 0 41768 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_457
timestamp 1644511149
transform 1 0 43148 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_464
timestamp 1644511149
transform 1 0 43792 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_471
timestamp 1644511149
transform 1 0 44436 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_496
timestamp 1644511149
transform 1 0 46736 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_512
timestamp 1644511149
transform 1 0 48208 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_520
timestamp 1644511149
transform 1 0 48944 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_536
timestamp 1644511149
transform 1 0 50416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_547
timestamp 1644511149
transform 1 0 51428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_555
timestamp 1644511149
transform 1 0 52164 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_565
timestamp 1644511149
transform 1 0 53084 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_588
timestamp 1644511149
transform 1 0 55200 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_598
timestamp 1644511149
transform 1 0 56120 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_606
timestamp 1644511149
transform 1 0 56856 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_614
timestamp 1644511149
transform 1 0 57592 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_620
timestamp 1644511149
transform 1 0 58144 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_624
timestamp 1644511149
transform 1 0 58512 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_259
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_276
timestamp 1644511149
transform 1 0 26496 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_288
timestamp 1644511149
transform 1 0 27600 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_296
timestamp 1644511149
transform 1 0 28336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_322
timestamp 1644511149
transform 1 0 30728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_342
timestamp 1644511149
transform 1 0 32568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1644511149
transform 1 0 33212 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_361
timestamp 1644511149
transform 1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_382
timestamp 1644511149
transform 1 0 36248 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_390
timestamp 1644511149
transform 1 0 36984 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_408
timestamp 1644511149
transform 1 0 38640 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_441
timestamp 1644511149
transform 1 0 41676 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_448
timestamp 1644511149
transform 1 0 42320 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_456
timestamp 1644511149
transform 1 0 43056 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_463
timestamp 1644511149
transform 1 0 43700 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_472
timestamp 1644511149
transform 1 0 44528 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_485
timestamp 1644511149
transform 1 0 45724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_497
timestamp 1644511149
transform 1 0 46828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_505
timestamp 1644511149
transform 1 0 47564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_521
timestamp 1644511149
transform 1 0 49036 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_529
timestamp 1644511149
transform 1 0 49772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_537
timestamp 1644511149
transform 1 0 50508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_548
timestamp 1644511149
transform 1 0 51520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_562
timestamp 1644511149
transform 1 0 52808 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_572
timestamp 1644511149
transform 1 0 53728 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_584
timestamp 1644511149
transform 1 0 54832 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_598
timestamp 1644511149
transform 1 0 56120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_610
timestamp 1644511149
transform 1 0 57224 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_622
timestamp 1644511149
transform 1 0 58328 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_274
timestamp 1644511149
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_284
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_296
timestamp 1644511149
transform 1 0 28336 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_304
timestamp 1644511149
transform 1 0 29072 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_316
timestamp 1644511149
transform 1 0 30176 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_328
timestamp 1644511149
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_342
timestamp 1644511149
transform 1 0 32568 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_354
timestamp 1644511149
transform 1 0 33672 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_358
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_375
timestamp 1644511149
transform 1 0 35604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 1644511149
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_409
timestamp 1644511149
transform 1 0 38732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_421
timestamp 1644511149
transform 1 0 39836 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_433
timestamp 1644511149
transform 1 0 40940 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_440
timestamp 1644511149
transform 1 0 41584 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_456
timestamp 1644511149
transform 1 0 43056 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_468
timestamp 1644511149
transform 1 0 44160 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_476
timestamp 1644511149
transform 1 0 44896 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_480
timestamp 1644511149
transform 1 0 45264 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_492
timestamp 1644511149
transform 1 0 46368 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_513
timestamp 1644511149
transform 1 0 48300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_522
timestamp 1644511149
transform 1 0 49128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_530
timestamp 1644511149
transform 1 0 49864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_536
timestamp 1644511149
transform 1 0 50416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_544
timestamp 1644511149
transform 1 0 51152 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_550
timestamp 1644511149
transform 1 0 51704 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_556
timestamp 1644511149
transform 1 0 52256 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_565
timestamp 1644511149
transform 1 0 53084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_572
timestamp 1644511149
transform 1 0 53728 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_584
timestamp 1644511149
transform 1 0 54832 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_592
timestamp 1644511149
transform 1 0 55568 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_603
timestamp 1644511149
transform 1 0 56580 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_610
timestamp 1644511149
transform 1 0 57224 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_269
timestamp 1644511149
transform 1 0 25852 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_282
timestamp 1644511149
transform 1 0 27048 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_318
timestamp 1644511149
transform 1 0 30360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_330
timestamp 1644511149
transform 1 0 31464 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_342
timestamp 1644511149
transform 1 0 32568 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 1644511149
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1644511149
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_385
timestamp 1644511149
transform 1 0 36524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_404
timestamp 1644511149
transform 1 0 38272 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_416
timestamp 1644511149
transform 1 0 39376 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_444
timestamp 1644511149
transform 1 0 41952 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_453
timestamp 1644511149
transform 1 0 42780 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_465
timestamp 1644511149
transform 1 0 43884 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_470
timestamp 1644511149
transform 1 0 44344 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_481
timestamp 1644511149
transform 1 0 45356 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_485
timestamp 1644511149
transform 1 0 45724 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_496
timestamp 1644511149
transform 1 0 46736 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_506
timestamp 1644511149
transform 1 0 47656 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_515
timestamp 1644511149
transform 1 0 48484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_527
timestamp 1644511149
transform 1 0 49588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_537
timestamp 1644511149
transform 1 0 50508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_546
timestamp 1644511149
transform 1 0 51336 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_554
timestamp 1644511149
transform 1 0 52072 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_566
timestamp 1644511149
transform 1 0 53176 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_572
timestamp 1644511149
transform 1 0 53728 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_577
timestamp 1644511149
transform 1 0 54188 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_584
timestamp 1644511149
transform 1 0 54832 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_596
timestamp 1644511149
transform 1 0 55936 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_621
timestamp 1644511149
transform 1 0 58236 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_245
timestamp 1644511149
transform 1 0 23644 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_253
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_262
timestamp 1644511149
transform 1 0 25208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1644511149
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_303
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_311
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_316
timestamp 1644511149
transform 1 0 30176 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_325
timestamp 1644511149
transform 1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1644511149
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_456
timestamp 1644511149
transform 1 0 43056 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_464
timestamp 1644511149
transform 1 0 43792 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_470
timestamp 1644511149
transform 1 0 44344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_478
timestamp 1644511149
transform 1 0 45080 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_510
timestamp 1644511149
transform 1 0 48024 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_518
timestamp 1644511149
transform 1 0 48760 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_524
timestamp 1644511149
transform 1 0 49312 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_532
timestamp 1644511149
transform 1 0 50048 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_542
timestamp 1644511149
transform 1 0 50968 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_549
timestamp 1644511149
transform 1 0 51612 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_557
timestamp 1644511149
transform 1 0 52348 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_579
timestamp 1644511149
transform 1 0 54372 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_587
timestamp 1644511149
transform 1 0 55108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_596
timestamp 1644511149
transform 1 0 55936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_604
timestamp 1644511149
transform 1 0 56672 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_611
timestamp 1644511149
transform 1 0 57316 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_620
timestamp 1644511149
transform 1 0 58144 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_624
timestamp 1644511149
transform 1 0 58512 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_259
timestamp 1644511149
transform 1 0 24932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_269
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_281
timestamp 1644511149
transform 1 0 26956 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_290
timestamp 1644511149
transform 1 0 27784 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_303
timestamp 1644511149
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_338
timestamp 1644511149
transform 1 0 32200 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_350
timestamp 1644511149
transform 1 0 33304 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1644511149
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_381
timestamp 1644511149
transform 1 0 36156 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_393
timestamp 1644511149
transform 1 0 37260 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_405
timestamp 1644511149
transform 1 0 38364 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_416
timestamp 1644511149
transform 1 0 39376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_425
timestamp 1644511149
transform 1 0 40204 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_435
timestamp 1644511149
transform 1 0 41124 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_447
timestamp 1644511149
transform 1 0 42228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_455
timestamp 1644511149
transform 1 0 42964 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_461
timestamp 1644511149
transform 1 0 43516 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_472
timestamp 1644511149
transform 1 0 44528 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_482
timestamp 1644511149
transform 1 0 45448 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_490
timestamp 1644511149
transform 1 0 46184 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_508
timestamp 1644511149
transform 1 0 47840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_517
timestamp 1644511149
transform 1 0 48668 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_527
timestamp 1644511149
transform 1 0 49588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_547
timestamp 1644511149
transform 1 0 51428 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_556
timestamp 1644511149
transform 1 0 52256 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_563
timestamp 1644511149
transform 1 0 52900 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_567
timestamp 1644511149
transform 1 0 53268 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_575
timestamp 1644511149
transform 1 0 54004 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_579
timestamp 1644511149
transform 1 0 54372 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_583
timestamp 1644511149
transform 1 0 54740 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_596
timestamp 1644511149
transform 1 0 55936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_621
timestamp 1644511149
transform 1 0 58236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_289
timestamp 1644511149
transform 1 0 27692 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_297
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_309
timestamp 1644511149
transform 1 0 29532 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_315
timestamp 1644511149
transform 1 0 30084 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_343
timestamp 1644511149
transform 1 0 32660 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_350
timestamp 1644511149
transform 1 0 33304 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_375
timestamp 1644511149
transform 1 0 35604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_387
timestamp 1644511149
transform 1 0 36708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_409
timestamp 1644511149
transform 1 0 38732 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_421
timestamp 1644511149
transform 1 0 39836 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_435
timestamp 1644511149
transform 1 0 41124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_444
timestamp 1644511149
transform 1 0 41952 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_472
timestamp 1644511149
transform 1 0 44528 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_482
timestamp 1644511149
transform 1 0 45448 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_489
timestamp 1644511149
transform 1 0 46092 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_500
timestamp 1644511149
transform 1 0 47104 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_515
timestamp 1644511149
transform 1 0 48484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_522
timestamp 1644511149
transform 1 0 49128 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_533
timestamp 1644511149
transform 1 0 50140 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_544
timestamp 1644511149
transform 1 0 51152 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_554
timestamp 1644511149
transform 1 0 52072 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_565
timestamp 1644511149
transform 1 0 53084 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_577
timestamp 1644511149
transform 1 0 54188 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_589
timestamp 1644511149
transform 1 0 55292 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_601
timestamp 1644511149
transform 1 0 56396 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_605
timestamp 1644511149
transform 1 0 56764 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_620
timestamp 1644511149
transform 1 0 58144 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_624
timestamp 1644511149
transform 1 0 58512 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_257
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_274
timestamp 1644511149
transform 1 0 26312 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_282
timestamp 1644511149
transform 1 0 27048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_287
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_293
timestamp 1644511149
transform 1 0 28060 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_341
timestamp 1644511149
transform 1 0 32476 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_353
timestamp 1644511149
transform 1 0 33580 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_361
timestamp 1644511149
transform 1 0 34316 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_381
timestamp 1644511149
transform 1 0 36156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_408
timestamp 1644511149
transform 1 0 38640 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_427
timestamp 1644511149
transform 1 0 40388 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_437
timestamp 1644511149
transform 1 0 41308 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_451
timestamp 1644511149
transform 1 0 42596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_471
timestamp 1644511149
transform 1 0 44436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_485
timestamp 1644511149
transform 1 0 45724 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_493
timestamp 1644511149
transform 1 0 46460 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_499
timestamp 1644511149
transform 1 0 47012 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_503
timestamp 1644511149
transform 1 0 47380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_515
timestamp 1644511149
transform 1 0 48484 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_548
timestamp 1644511149
transform 1 0 51520 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_554
timestamp 1644511149
transform 1 0 52072 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_562
timestamp 1644511149
transform 1 0 52808 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_597
timestamp 1644511149
transform 1 0 56028 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_602
timestamp 1644511149
transform 1 0 56488 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_611
timestamp 1644511149
transform 1 0 57316 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_623
timestamp 1644511149
transform 1 0 58420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_257
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_287
timestamp 1644511149
transform 1 0 27508 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_307
timestamp 1644511149
transform 1 0 29348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_319
timestamp 1644511149
transform 1 0 30452 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1644511149
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_345
timestamp 1644511149
transform 1 0 32844 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_357
timestamp 1644511149
transform 1 0 33948 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_366
timestamp 1644511149
transform 1 0 34776 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_409
timestamp 1644511149
transform 1 0 38732 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_421
timestamp 1644511149
transform 1 0 39836 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_432
timestamp 1644511149
transform 1 0 40848 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_442
timestamp 1644511149
transform 1 0 41768 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_456
timestamp 1644511149
transform 1 0 43056 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_465
timestamp 1644511149
transform 1 0 43884 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_474
timestamp 1644511149
transform 1 0 44712 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_482
timestamp 1644511149
transform 1 0 45448 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_494
timestamp 1644511149
transform 1 0 46552 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_502
timestamp 1644511149
transform 1 0 47288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_509
timestamp 1644511149
transform 1 0 47932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_525
timestamp 1644511149
transform 1 0 49404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_534
timestamp 1644511149
transform 1 0 50232 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_542
timestamp 1644511149
transform 1 0 50968 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_546
timestamp 1644511149
transform 1 0 51336 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_551
timestamp 1644511149
transform 1 0 51796 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_593
timestamp 1644511149
transform 1 0 55660 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_604
timestamp 1644511149
transform 1 0 56672 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1644511149
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_279
timestamp 1644511149
transform 1 0 26772 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_303
timestamp 1644511149
transform 1 0 28980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_319
timestamp 1644511149
transform 1 0 30452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_323
timestamp 1644511149
transform 1 0 30820 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_340
timestamp 1644511149
transform 1 0 32384 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_348
timestamp 1644511149
transform 1 0 33120 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_356
timestamp 1644511149
transform 1 0 33856 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_372
timestamp 1644511149
transform 1 0 35328 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_379
timestamp 1644511149
transform 1 0 35972 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_391
timestamp 1644511149
transform 1 0 37076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_415
timestamp 1644511149
transform 1 0 39284 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_453
timestamp 1644511149
transform 1 0 42780 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_462
timestamp 1644511149
transform 1 0 43608 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_470
timestamp 1644511149
transform 1 0 44344 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_492
timestamp 1644511149
transform 1 0 46368 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_506
timestamp 1644511149
transform 1 0 47656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_517
timestamp 1644511149
transform 1 0 48668 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_529
timestamp 1644511149
transform 1 0 49772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_553
timestamp 1644511149
transform 1 0 51980 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_562
timestamp 1644511149
transform 1 0 52808 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_573
timestamp 1644511149
transform 1 0 53820 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_585
timestamp 1644511149
transform 1 0 54924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_602
timestamp 1644511149
transform 1 0 56488 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_611
timestamp 1644511149
transform 1 0 57316 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1644511149
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_232
timestamp 1644511149
transform 1 0 22448 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_240
timestamp 1644511149
transform 1 0 23184 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_252
timestamp 1644511149
transform 1 0 24288 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_264
timestamp 1644511149
transform 1 0 25392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1644511149
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_301
timestamp 1644511149
transform 1 0 28796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_311
timestamp 1644511149
transform 1 0 29716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_323
timestamp 1644511149
transform 1 0 30820 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_354
timestamp 1644511149
transform 1 0 33672 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_365
timestamp 1644511149
transform 1 0 34684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_376
timestamp 1644511149
transform 1 0 35696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_380
timestamp 1644511149
transform 1 0 36064 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1644511149
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_400
timestamp 1644511149
transform 1 0 37904 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_412
timestamp 1644511149
transform 1 0 39008 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_424
timestamp 1644511149
transform 1 0 40112 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_432
timestamp 1644511149
transform 1 0 40848 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_437
timestamp 1644511149
transform 1 0 41308 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_445
timestamp 1644511149
transform 1 0 42044 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_469
timestamp 1644511149
transform 1 0 44252 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_476
timestamp 1644511149
transform 1 0 44896 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_488
timestamp 1644511149
transform 1 0 46000 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_500
timestamp 1644511149
transform 1 0 47104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_510
timestamp 1644511149
transform 1 0 48024 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_522
timestamp 1644511149
transform 1 0 49128 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_528
timestamp 1644511149
transform 1 0 49680 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_534
timestamp 1644511149
transform 1 0 50232 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_580
timestamp 1644511149
transform 1 0 54464 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_591
timestamp 1644511149
transform 1 0 55476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_602
timestamp 1644511149
transform 1 0 56488 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_612
timestamp 1644511149
transform 1 0 57408 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_620
timestamp 1644511149
transform 1 0 58144 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_624
timestamp 1644511149
transform 1 0 58512 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_205
timestamp 1644511149
transform 1 0 19964 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_214
timestamp 1644511149
transform 1 0 20792 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_236
timestamp 1644511149
transform 1 0 22816 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1644511149
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_286
timestamp 1644511149
transform 1 0 27416 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_292
timestamp 1644511149
transform 1 0 27968 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_297
timestamp 1644511149
transform 1 0 28428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1644511149
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_338
timestamp 1644511149
transform 1 0 32200 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_375
timestamp 1644511149
transform 1 0 35604 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_383
timestamp 1644511149
transform 1 0 36340 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1644511149
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_406
timestamp 1644511149
transform 1 0 38456 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_418
timestamp 1644511149
transform 1 0 39560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_425
timestamp 1644511149
transform 1 0 40204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_436
timestamp 1644511149
transform 1 0 41216 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_448
timestamp 1644511149
transform 1 0 42320 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_454
timestamp 1644511149
transform 1 0 42872 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_464
timestamp 1644511149
transform 1 0 43792 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_483
timestamp 1644511149
transform 1 0 45540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_491
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_504
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_518
timestamp 1644511149
transform 1 0 48760 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_526
timestamp 1644511149
transform 1 0 49496 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_540
timestamp 1644511149
transform 1 0 50784 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_552
timestamp 1644511149
transform 1 0 51888 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_564
timestamp 1644511149
transform 1 0 52992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_576
timestamp 1644511149
transform 1 0 54096 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_597
timestamp 1644511149
transform 1 0 56028 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_612
timestamp 1644511149
transform 1 0 57408 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_620
timestamp 1644511149
transform 1 0 58144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_624
timestamp 1644511149
transform 1 0 58512 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_201
timestamp 1644511149
transform 1 0 19596 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_211
timestamp 1644511149
transform 1 0 20516 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_215
timestamp 1644511149
transform 1 0 20884 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_235
timestamp 1644511149
transform 1 0 22724 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_246
timestamp 1644511149
transform 1 0 23736 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_259
timestamp 1644511149
transform 1 0 24932 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_268
timestamp 1644511149
transform 1 0 25760 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_275
timestamp 1644511149
transform 1 0 26404 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_309
timestamp 1644511149
transform 1 0 29532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_321
timestamp 1644511149
transform 1 0 30636 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1644511149
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_345
timestamp 1644511149
transform 1 0 32844 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_359
timestamp 1644511149
transform 1 0 34132 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_388
timestamp 1644511149
transform 1 0 36800 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_403
timestamp 1644511149
transform 1 0 38180 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_414
timestamp 1644511149
transform 1 0 39192 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_435
timestamp 1644511149
transform 1 0 41124 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_443
timestamp 1644511149
transform 1 0 41860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_454
timestamp 1644511149
transform 1 0 42872 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_467
timestamp 1644511149
transform 1 0 44068 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_477
timestamp 1644511149
transform 1 0 44988 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_494
timestamp 1644511149
transform 1 0 46552 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_502
timestamp 1644511149
transform 1 0 47288 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_510
timestamp 1644511149
transform 1 0 48024 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_523
timestamp 1644511149
transform 1 0 49220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_533
timestamp 1644511149
transform 1 0 50140 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_547
timestamp 1644511149
transform 1 0 51428 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_556
timestamp 1644511149
transform 1 0 52256 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_570
timestamp 1644511149
transform 1 0 53544 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_582
timestamp 1644511149
transform 1 0 54648 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_594
timestamp 1644511149
transform 1 0 55752 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_602
timestamp 1644511149
transform 1 0 56488 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_610
timestamp 1644511149
transform 1 0 57224 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_213
timestamp 1644511149
transform 1 0 20700 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_231
timestamp 1644511149
transform 1 0 22356 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_241
timestamp 1644511149
transform 1 0 23276 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1644511149
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_262
timestamp 1644511149
transform 1 0 25208 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_274
timestamp 1644511149
transform 1 0 26312 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_279
timestamp 1644511149
transform 1 0 26772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_291
timestamp 1644511149
transform 1 0 27876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_303
timestamp 1644511149
transform 1 0 28980 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_317
timestamp 1644511149
transform 1 0 30268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_326
timestamp 1644511149
transform 1 0 31096 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_334
timestamp 1644511149
transform 1 0 31832 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_350
timestamp 1644511149
transform 1 0 33304 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_372
timestamp 1644511149
transform 1 0 35328 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_379
timestamp 1644511149
transform 1 0 35972 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_383
timestamp 1644511149
transform 1 0 36340 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_391
timestamp 1644511149
transform 1 0 37076 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_402
timestamp 1644511149
transform 1 0 38088 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_443
timestamp 1644511149
transform 1 0 41860 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_455
timestamp 1644511149
transform 1 0 42964 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_466
timestamp 1644511149
transform 1 0 43976 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_474
timestamp 1644511149
transform 1 0 44712 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_487
timestamp 1644511149
transform 1 0 45908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_499
timestamp 1644511149
transform 1 0 47012 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_507
timestamp 1644511149
transform 1 0 47748 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_516
timestamp 1644511149
transform 1 0 48576 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_524
timestamp 1644511149
transform 1 0 49312 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_528
timestamp 1644511149
transform 1 0 49680 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_543
timestamp 1644511149
transform 1 0 51060 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_552
timestamp 1644511149
transform 1 0 51888 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_565
timestamp 1644511149
transform 1 0 53084 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_573
timestamp 1644511149
transform 1 0 53820 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_585
timestamp 1644511149
transform 1 0 54924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_597
timestamp 1644511149
transform 1 0 56028 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_621
timestamp 1644511149
transform 1 0 58236 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_11
timestamp 1644511149
transform 1 0 2116 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_33
timestamp 1644511149
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1644511149
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1644511149
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_211
timestamp 1644511149
transform 1 0 20516 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 1644511149
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_231
timestamp 1644511149
transform 1 0 22356 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_239
timestamp 1644511149
transform 1 0 23092 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_245
timestamp 1644511149
transform 1 0 23644 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_250
timestamp 1644511149
transform 1 0 24104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_254
timestamp 1644511149
transform 1 0 24472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_265
timestamp 1644511149
transform 1 0 25484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_277
timestamp 1644511149
transform 1 0 26588 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_289
timestamp 1644511149
transform 1 0 27692 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_304
timestamp 1644511149
transform 1 0 29072 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_316
timestamp 1644511149
transform 1 0 30176 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_325
timestamp 1644511149
transform 1 0 31004 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1644511149
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_348
timestamp 1644511149
transform 1 0 33120 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_355
timestamp 1644511149
transform 1 0 33764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_368
timestamp 1644511149
transform 1 0 34960 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_375
timestamp 1644511149
transform 1 0 35604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_387
timestamp 1644511149
transform 1 0 36708 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_400
timestamp 1644511149
transform 1 0 37904 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_408
timestamp 1644511149
transform 1 0 38640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_416
timestamp 1644511149
transform 1 0 39376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_425
timestamp 1644511149
transform 1 0 40204 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_434
timestamp 1644511149
transform 1 0 41032 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_442
timestamp 1644511149
transform 1 0 41768 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_457
timestamp 1644511149
transform 1 0 43148 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_467
timestamp 1644511149
transform 1 0 44068 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_480
timestamp 1644511149
transform 1 0 45264 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_492
timestamp 1644511149
transform 1 0 46368 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_511
timestamp 1644511149
transform 1 0 48116 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_516
timestamp 1644511149
transform 1 0 48576 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_527
timestamp 1644511149
transform 1 0 49588 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_535
timestamp 1644511149
transform 1 0 50324 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_549
timestamp 1644511149
transform 1 0 51612 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_556
timestamp 1644511149
transform 1 0 52256 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_570
timestamp 1644511149
transform 1 0 53544 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_582
timestamp 1644511149
transform 1 0 54648 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_594
timestamp 1644511149
transform 1 0 55752 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_606
timestamp 1644511149
transform 1 0 56856 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_614
timestamp 1644511149
transform 1 0 57592 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_620
timestamp 1644511149
transform 1 0 58144 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_624
timestamp 1644511149
transform 1 0 58512 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1644511149
transform 1 0 4048 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1644511149
transform 1 0 5152 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_56
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_68
timestamp 1644511149
transform 1 0 7360 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1644511149
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_218
timestamp 1644511149
transform 1 0 21160 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_230
timestamp 1644511149
transform 1 0 22264 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_234
timestamp 1644511149
transform 1 0 22632 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_238
timestamp 1644511149
transform 1 0 23000 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1644511149
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_261
timestamp 1644511149
transform 1 0 25116 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_269
timestamp 1644511149
transform 1 0 25852 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_281
timestamp 1644511149
transform 1 0 26956 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_287
timestamp 1644511149
transform 1 0 27508 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_304
timestamp 1644511149
transform 1 0 29072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_316
timestamp 1644511149
transform 1 0 30176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_324
timestamp 1644511149
transform 1 0 30912 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_332
timestamp 1644511149
transform 1 0 31648 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_341
timestamp 1644511149
transform 1 0 32476 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_353
timestamp 1644511149
transform 1 0 33580 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1644511149
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_372
timestamp 1644511149
transform 1 0 35328 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_384
timestamp 1644511149
transform 1 0 36432 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_396
timestamp 1644511149
transform 1 0 37536 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_408
timestamp 1644511149
transform 1 0 38640 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_427
timestamp 1644511149
transform 1 0 40388 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_435
timestamp 1644511149
transform 1 0 41124 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_447
timestamp 1644511149
transform 1 0 42228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_459
timestamp 1644511149
transform 1 0 43332 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_472
timestamp 1644511149
transform 1 0 44528 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_485
timestamp 1644511149
transform 1 0 45724 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_497
timestamp 1644511149
transform 1 0 46828 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_509
timestamp 1644511149
transform 1 0 47932 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_513
timestamp 1644511149
transform 1 0 48300 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_521
timestamp 1644511149
transform 1 0 49036 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_529
timestamp 1644511149
transform 1 0 49772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_537
timestamp 1644511149
transform 1 0 50508 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_551
timestamp 1644511149
transform 1 0 51796 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_563
timestamp 1644511149
transform 1 0 52900 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_575
timestamp 1644511149
transform 1 0 54004 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_584
timestamp 1644511149
transform 1 0 54832 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_595
timestamp 1644511149
transform 1 0 55844 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_599
timestamp 1644511149
transform 1 0 56212 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_606
timestamp 1644511149
transform 1 0 56856 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_613
timestamp 1644511149
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_11
timestamp 1644511149
transform 1 0 2116 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_233
timestamp 1644511149
transform 1 0 22540 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_241
timestamp 1644511149
transform 1 0 23276 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_269
timestamp 1644511149
transform 1 0 25852 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 1644511149
transform 1 0 26496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_289
timestamp 1644511149
transform 1 0 27692 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_303
timestamp 1644511149
transform 1 0 28980 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_311
timestamp 1644511149
transform 1 0 29716 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_326
timestamp 1644511149
transform 1 0 31096 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 1644511149
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_341
timestamp 1644511149
transform 1 0 32476 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_353
timestamp 1644511149
transform 1 0 33580 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_369
timestamp 1644511149
transform 1 0 35052 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_381
timestamp 1644511149
transform 1 0 36156 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_389
timestamp 1644511149
transform 1 0 36892 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_401
timestamp 1644511149
transform 1 0 37996 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_408
timestamp 1644511149
transform 1 0 38640 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_416
timestamp 1644511149
transform 1 0 39376 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_421
timestamp 1644511149
transform 1 0 39836 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_434
timestamp 1644511149
transform 1 0 41032 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_443
timestamp 1644511149
transform 1 0 41860 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_471
timestamp 1644511149
transform 1 0 44436 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_475
timestamp 1644511149
transform 1 0 44804 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_483
timestamp 1644511149
transform 1 0 45540 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_495
timestamp 1644511149
transform 1 0 46644 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_500
timestamp 1644511149
transform 1 0 47104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_505
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_513
timestamp 1644511149
transform 1 0 48300 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_521
timestamp 1644511149
transform 1 0 49036 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_526
timestamp 1644511149
transform 1 0 49496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_533
timestamp 1644511149
transform 1 0 50140 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_537
timestamp 1644511149
transform 1 0 50508 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_541
timestamp 1644511149
transform 1 0 50876 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_552
timestamp 1644511149
transform 1 0 51888 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_568
timestamp 1644511149
transform 1 0 53360 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_577
timestamp 1644511149
transform 1 0 54188 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_588
timestamp 1644511149
transform 1 0 55200 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_603
timestamp 1644511149
transform 1 0 56580 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1644511149
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_621
timestamp 1644511149
transform 1 0 58236 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_215
timestamp 1644511149
transform 1 0 20884 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_220
timestamp 1644511149
transform 1 0 21344 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_227
timestamp 1644511149
transform 1 0 21988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_243
timestamp 1644511149
transform 1 0 23460 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_259
timestamp 1644511149
transform 1 0 24932 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_268
timestamp 1644511149
transform 1 0 25760 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_280
timestamp 1644511149
transform 1 0 26864 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_286
timestamp 1644511149
transform 1 0 27416 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_290
timestamp 1644511149
transform 1 0 27784 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1644511149
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_322
timestamp 1644511149
transform 1 0 30728 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_331
timestamp 1644511149
transform 1 0 31556 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_353
timestamp 1644511149
transform 1 0 33580 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_361
timestamp 1644511149
transform 1 0 34316 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_371
timestamp 1644511149
transform 1 0 35236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_383
timestamp 1644511149
transform 1 0 36340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_393
timestamp 1644511149
transform 1 0 37260 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_405
timestamp 1644511149
transform 1 0 38364 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_416
timestamp 1644511149
transform 1 0 39376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_429
timestamp 1644511149
transform 1 0 40572 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_442
timestamp 1644511149
transform 1 0 41768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_449
timestamp 1644511149
transform 1 0 42412 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_497
timestamp 1644511149
transform 1 0 46828 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_509
timestamp 1644511149
transform 1 0 47932 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_516
timestamp 1644511149
transform 1 0 48576 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_528
timestamp 1644511149
transform 1 0 49680 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_538
timestamp 1644511149
transform 1 0 50600 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_553
timestamp 1644511149
transform 1 0 51980 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_561
timestamp 1644511149
transform 1 0 52716 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_573
timestamp 1644511149
transform 1 0 53820 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_585
timestamp 1644511149
transform 1 0 54924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_595
timestamp 1644511149
transform 1 0 55844 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_599
timestamp 1644511149
transform 1 0 56212 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_605
timestamp 1644511149
transform 1 0 56764 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_612
timestamp 1644511149
transform 1 0 57408 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_624
timestamp 1644511149
transform 1 0 58512 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_209
timestamp 1644511149
transform 1 0 20332 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_230
timestamp 1644511149
transform 1 0 22264 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_242
timestamp 1644511149
transform 1 0 23368 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_251
timestamp 1644511149
transform 1 0 24196 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_259
timestamp 1644511149
transform 1 0 24932 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_271
timestamp 1644511149
transform 1 0 26036 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_287
timestamp 1644511149
transform 1 0 27508 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_300
timestamp 1644511149
transform 1 0 28704 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_308
timestamp 1644511149
transform 1 0 29440 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_313
timestamp 1644511149
transform 1 0 29900 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_327
timestamp 1644511149
transform 1 0 31188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_344
timestamp 1644511149
transform 1 0 32752 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_353
timestamp 1644511149
transform 1 0 33580 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_360
timestamp 1644511149
transform 1 0 34224 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_372
timestamp 1644511149
transform 1 0 35328 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_384
timestamp 1644511149
transform 1 0 36432 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_406
timestamp 1644511149
transform 1 0 38456 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_415
timestamp 1644511149
transform 1 0 39284 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_424
timestamp 1644511149
transform 1 0 40112 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_433
timestamp 1644511149
transform 1 0 40940 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_71_442
timestamp 1644511149
transform 1 0 41768 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_458
timestamp 1644511149
transform 1 0 43240 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_470
timestamp 1644511149
transform 1 0 44344 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_482
timestamp 1644511149
transform 1 0 45448 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_494
timestamp 1644511149
transform 1 0 46552 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1644511149
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_515
timestamp 1644511149
transform 1 0 48484 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_524
timestamp 1644511149
transform 1 0 49312 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_538
timestamp 1644511149
transform 1 0 50600 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_549
timestamp 1644511149
transform 1 0 51612 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_556
timestamp 1644511149
transform 1 0 52256 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_561
timestamp 1644511149
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_573
timestamp 1644511149
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_585
timestamp 1644511149
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_597
timestamp 1644511149
transform 1 0 56028 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_602
timestamp 1644511149
transform 1 0 56488 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_611
timestamp 1644511149
transform 1 0 57316 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1644511149
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1644511149
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_203
timestamp 1644511149
transform 1 0 19780 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_215
timestamp 1644511149
transform 1 0 20884 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_227
timestamp 1644511149
transform 1 0 21988 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_237
timestamp 1644511149
transform 1 0 22908 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_243
timestamp 1644511149
transform 1 0 23460 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1644511149
transform 1 0 23920 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_261
timestamp 1644511149
transform 1 0 25116 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_273
timestamp 1644511149
transform 1 0 26220 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_285
timestamp 1644511149
transform 1 0 27324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_294
timestamp 1644511149
transform 1 0 28152 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1644511149
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_331
timestamp 1644511149
transform 1 0 31556 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_343
timestamp 1644511149
transform 1 0 32660 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_353
timestamp 1644511149
transform 1 0 33580 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1644511149
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_397
timestamp 1644511149
transform 1 0 37628 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_409
timestamp 1644511149
transform 1 0 38732 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_417
timestamp 1644511149
transform 1 0 39468 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_452
timestamp 1644511149
transform 1 0 42688 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_464
timestamp 1644511149
transform 1 0 43792 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_482
timestamp 1644511149
transform 1 0 45448 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_494
timestamp 1644511149
transform 1 0 46552 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_502
timestamp 1644511149
transform 1 0 47288 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_510
timestamp 1644511149
transform 1 0 48024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_518
timestamp 1644511149
transform 1 0 48760 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_530
timestamp 1644511149
transform 1 0 49864 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_533
timestamp 1644511149
transform 1 0 50140 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_540
timestamp 1644511149
transform 1 0 50784 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_547
timestamp 1644511149
transform 1 0 51428 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_559
timestamp 1644511149
transform 1 0 52532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_571
timestamp 1644511149
transform 1 0 53636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_583
timestamp 1644511149
transform 1 0 54740 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1644511149
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_589
timestamp 1644511149
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_601
timestamp 1644511149
transform 1 0 56396 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_608
timestamp 1644511149
transform 1 0 57040 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_620
timestamp 1644511149
transform 1 0 58144 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_624
timestamp 1644511149
transform 1 0 58512 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_199
timestamp 1644511149
transform 1 0 19412 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_216
timestamp 1644511149
transform 1 0 20976 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_232
timestamp 1644511149
transform 1 0 22448 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_244
timestamp 1644511149
transform 1 0 23552 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_263
timestamp 1644511149
transform 1 0 25300 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_267
timestamp 1644511149
transform 1 0 25668 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1644511149
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_291
timestamp 1644511149
transform 1 0 27876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_315
timestamp 1644511149
transform 1 0 30084 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_322
timestamp 1644511149
transform 1 0 30728 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_326
timestamp 1644511149
transform 1 0 31096 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_330
timestamp 1644511149
transform 1 0 31464 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_344
timestamp 1644511149
transform 1 0 32752 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_356
timestamp 1644511149
transform 1 0 33856 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_376
timestamp 1644511149
transform 1 0 35696 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_388
timestamp 1644511149
transform 1 0 36800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_401
timestamp 1644511149
transform 1 0 37996 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_409
timestamp 1644511149
transform 1 0 38732 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_418
timestamp 1644511149
transform 1 0 39560 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_426
timestamp 1644511149
transform 1 0 40296 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_433
timestamp 1644511149
transform 1 0 40940 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_439
timestamp 1644511149
transform 1 0 41492 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_444
timestamp 1644511149
transform 1 0 41952 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_454
timestamp 1644511149
transform 1 0 42872 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_505
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_511
timestamp 1644511149
transform 1 0 48116 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_518
timestamp 1644511149
transform 1 0 48760 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_530
timestamp 1644511149
transform 1 0 49864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_534
timestamp 1644511149
transform 1 0 50232 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_546
timestamp 1644511149
transform 1 0 51336 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1644511149
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1644511149
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_561
timestamp 1644511149
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_573
timestamp 1644511149
transform 1 0 53820 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_581
timestamp 1644511149
transform 1 0 54556 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_591
timestamp 1644511149
transform 1 0 55476 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_603
timestamp 1644511149
transform 1 0 56580 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1644511149
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1644511149
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_620
timestamp 1644511149
transform 1 0 58144 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_624
timestamp 1644511149
transform 1 0 58512 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_205
timestamp 1644511149
transform 1 0 19964 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_213
timestamp 1644511149
transform 1 0 20700 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_217
timestamp 1644511149
transform 1 0 21068 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_234
timestamp 1644511149
transform 1 0 22632 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_240
timestamp 1644511149
transform 1 0 23184 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_248
timestamp 1644511149
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_257
timestamp 1644511149
transform 1 0 24748 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_279
timestamp 1644511149
transform 1 0 26772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_287
timestamp 1644511149
transform 1 0 27508 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_296
timestamp 1644511149
transform 1 0 28336 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_312
timestamp 1644511149
transform 1 0 29808 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_329
timestamp 1644511149
transform 1 0 31372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_336
timestamp 1644511149
transform 1 0 32016 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_344
timestamp 1644511149
transform 1 0 32752 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_356
timestamp 1644511149
transform 1 0 33856 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_381
timestamp 1644511149
transform 1 0 36156 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_400
timestamp 1644511149
transform 1 0 37904 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_411
timestamp 1644511149
transform 1 0 38916 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_454
timestamp 1644511149
transform 1 0 42872 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_466
timestamp 1644511149
transform 1 0 43976 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_474
timestamp 1644511149
transform 1 0 44712 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_486
timestamp 1644511149
transform 1 0 45816 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_490
timestamp 1644511149
transform 1 0 46184 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_496
timestamp 1644511149
transform 1 0 46736 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_503
timestamp 1644511149
transform 1 0 47380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_514
timestamp 1644511149
transform 1 0 48392 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_526
timestamp 1644511149
transform 1 0 49496 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_533
timestamp 1644511149
transform 1 0 50140 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_541
timestamp 1644511149
transform 1 0 50876 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_548
timestamp 1644511149
transform 1 0 51520 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_556
timestamp 1644511149
transform 1 0 52256 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_566
timestamp 1644511149
transform 1 0 53176 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_574
timestamp 1644511149
transform 1 0 53912 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_580
timestamp 1644511149
transform 1 0 54464 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_593
timestamp 1644511149
transform 1 0 55660 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_599
timestamp 1644511149
transform 1 0 56212 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_621
timestamp 1644511149
transform 1 0 58236 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_235
timestamp 1644511149
transform 1 0 22724 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_243
timestamp 1644511149
transform 1 0 23460 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_247
timestamp 1644511149
transform 1 0 23828 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_255
timestamp 1644511149
transform 1 0 24564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_266
timestamp 1644511149
transform 1 0 25576 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1644511149
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_365
timestamp 1644511149
transform 1 0 34684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_375
timestamp 1644511149
transform 1 0 35604 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_388
timestamp 1644511149
transform 1 0 36800 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_409
timestamp 1644511149
transform 1 0 38732 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_421
timestamp 1644511149
transform 1 0 39836 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_442
timestamp 1644511149
transform 1 0 41768 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_458
timestamp 1644511149
transform 1 0 43240 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_466
timestamp 1644511149
transform 1 0 43976 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_476
timestamp 1644511149
transform 1 0 44896 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_489
timestamp 1644511149
transform 1 0 46092 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_499
timestamp 1644511149
transform 1 0 47012 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1644511149
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_509
timestamp 1644511149
transform 1 0 47932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_531
timestamp 1644511149
transform 1 0 49956 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_543
timestamp 1644511149
transform 1 0 51060 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_551
timestamp 1644511149
transform 1 0 51796 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1644511149
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_571
timestamp 1644511149
transform 1 0 53636 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_75_580
timestamp 1644511149
transform 1 0 54464 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_586
timestamp 1644511149
transform 1 0 55016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_593
timestamp 1644511149
transform 1 0 55660 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_610
timestamp 1644511149
transform 1 0 57224 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_620
timestamp 1644511149
transform 1 0 58144 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_624
timestamp 1644511149
transform 1 0 58512 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_295
timestamp 1644511149
transform 1 0 28244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_312
timestamp 1644511149
transform 1 0 29808 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_324
timestamp 1644511149
transform 1 0 30912 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_342
timestamp 1644511149
transform 1 0 32568 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_354
timestamp 1644511149
transform 1 0 33672 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1644511149
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_373
timestamp 1644511149
transform 1 0 35420 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_384
timestamp 1644511149
transform 1 0 36432 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_396
timestamp 1644511149
transform 1 0 37536 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_405
timestamp 1644511149
transform 1 0 38364 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_416
timestamp 1644511149
transform 1 0 39376 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_428
timestamp 1644511149
transform 1 0 40480 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_434
timestamp 1644511149
transform 1 0 41032 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_442
timestamp 1644511149
transform 1 0 41768 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_472
timestamp 1644511149
transform 1 0 44528 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_485
timestamp 1644511149
transform 1 0 45724 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_497
timestamp 1644511149
transform 1 0 46828 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_508
timestamp 1644511149
transform 1 0 47840 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_515
timestamp 1644511149
transform 1 0 48484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_527
timestamp 1644511149
transform 1 0 49588 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1644511149
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_541
timestamp 1644511149
transform 1 0 50876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_553
timestamp 1644511149
transform 1 0 51980 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_561
timestamp 1644511149
transform 1 0 52716 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_569
timestamp 1644511149
transform 1 0 53452 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_575
timestamp 1644511149
transform 1 0 54004 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_584
timestamp 1644511149
transform 1 0 54832 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_594
timestamp 1644511149
transform 1 0 55752 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_621
timestamp 1644511149
transform 1 0 58236 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_199
timestamp 1644511149
transform 1 0 19412 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_203
timestamp 1644511149
transform 1 0 19780 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_215
timestamp 1644511149
transform 1 0 20884 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_253
timestamp 1644511149
transform 1 0 24380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_309
timestamp 1644511149
transform 1 0 29532 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_321
timestamp 1644511149
transform 1 0 30636 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_333
timestamp 1644511149
transform 1 0 31740 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_345
timestamp 1644511149
transform 1 0 32844 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_351
timestamp 1644511149
transform 1 0 33396 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_368
timestamp 1644511149
transform 1 0 34960 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_380
timestamp 1644511149
transform 1 0 36064 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_422
timestamp 1644511149
transform 1 0 39928 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_434
timestamp 1644511149
transform 1 0 41032 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_440
timestamp 1644511149
transform 1 0 41584 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_456
timestamp 1644511149
transform 1 0 43056 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_464
timestamp 1644511149
transform 1 0 43792 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_472
timestamp 1644511149
transform 1 0 44528 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_478
timestamp 1644511149
transform 1 0 45080 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1644511149
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_505
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_513
timestamp 1644511149
transform 1 0 48300 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_521
timestamp 1644511149
transform 1 0 49036 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_525
timestamp 1644511149
transform 1 0 49404 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_531
timestamp 1644511149
transform 1 0 49956 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_535
timestamp 1644511149
transform 1 0 50324 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_539
timestamp 1644511149
transform 1 0 50692 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_545
timestamp 1644511149
transform 1 0 51244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_556
timestamp 1644511149
transform 1 0 52256 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_566
timestamp 1644511149
transform 1 0 53176 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_573
timestamp 1644511149
transform 1 0 53820 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_579
timestamp 1644511149
transform 1 0 54372 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_584
timestamp 1644511149
transform 1 0 54832 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_596
timestamp 1644511149
transform 1 0 55936 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_606
timestamp 1644511149
transform 1 0 56856 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_614
timestamp 1644511149
transform 1 0 57592 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_620
timestamp 1644511149
transform 1 0 58144 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_624
timestamp 1644511149
transform 1 0 58512 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_200
timestamp 1644511149
transform 1 0 19504 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_212
timestamp 1644511149
transform 1 0 20608 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_224
timestamp 1644511149
transform 1 0 21712 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_236
timestamp 1644511149
transform 1 0 22816 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1644511149
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_261
timestamp 1644511149
transform 1 0 25116 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_270
timestamp 1644511149
transform 1 0 25944 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_282
timestamp 1644511149
transform 1 0 27048 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_288
timestamp 1644511149
transform 1 0 27600 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1644511149
transform 1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_314
timestamp 1644511149
transform 1 0 29992 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_338
timestamp 1644511149
transform 1 0 32200 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_350
timestamp 1644511149
transform 1 0 33304 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_362
timestamp 1644511149
transform 1 0 34408 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_381
timestamp 1644511149
transform 1 0 36156 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_398
timestamp 1644511149
transform 1 0 37720 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_409
timestamp 1644511149
transform 1 0 38732 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_416
timestamp 1644511149
transform 1 0 39376 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_425
timestamp 1644511149
transform 1 0 40204 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_434
timestamp 1644511149
transform 1 0 41032 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_442
timestamp 1644511149
transform 1 0 41768 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_450
timestamp 1644511149
transform 1 0 42504 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_459
timestamp 1644511149
transform 1 0 43332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_471
timestamp 1644511149
transform 1 0 44436 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_485
timestamp 1644511149
transform 1 0 45724 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_499
timestamp 1644511149
transform 1 0 47012 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_520
timestamp 1644511149
transform 1 0 48944 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_528
timestamp 1644511149
transform 1 0 49680 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_533
timestamp 1644511149
transform 1 0 50140 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_543
timestamp 1644511149
transform 1 0 51060 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_555
timestamp 1644511149
transform 1 0 52164 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_565
timestamp 1644511149
transform 1 0 53084 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_572
timestamp 1644511149
transform 1 0 53728 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_584
timestamp 1644511149
transform 1 0 54832 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_596
timestamp 1644511149
transform 1 0 55936 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_621
timestamp 1644511149
transform 1 0 58236 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_209
timestamp 1644511149
transform 1 0 20332 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 1644511149
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_247
timestamp 1644511149
transform 1 0 23828 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_257
timestamp 1644511149
transform 1 0 24748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_267
timestamp 1644511149
transform 1 0 25668 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_274
timestamp 1644511149
transform 1 0 26312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_290
timestamp 1644511149
transform 1 0 27784 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_310
timestamp 1644511149
transform 1 0 29624 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_318
timestamp 1644511149
transform 1 0 30360 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_330
timestamp 1644511149
transform 1 0 31464 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_79_353
timestamp 1644511149
transform 1 0 33580 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_364
timestamp 1644511149
transform 1 0 34592 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_377
timestamp 1644511149
transform 1 0 35788 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_383
timestamp 1644511149
transform 1 0 36340 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_401
timestamp 1644511149
transform 1 0 37996 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_412
timestamp 1644511149
transform 1 0 39008 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_424
timestamp 1644511149
transform 1 0 40112 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_433
timestamp 1644511149
transform 1 0 40940 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_444
timestamp 1644511149
transform 1 0 41952 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_458
timestamp 1644511149
transform 1 0 43240 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_470
timestamp 1644511149
transform 1 0 44344 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_482
timestamp 1644511149
transform 1 0 45448 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_489
timestamp 1644511149
transform 1 0 46092 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_495
timestamp 1644511149
transform 1 0 46644 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_499
timestamp 1644511149
transform 1 0 47012 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1644511149
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1644511149
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_526
timestamp 1644511149
transform 1 0 49496 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_538
timestamp 1644511149
transform 1 0 50600 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_544
timestamp 1644511149
transform 1 0 51152 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_552
timestamp 1644511149
transform 1 0 51888 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_561
timestamp 1644511149
transform 1 0 52716 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_569
timestamp 1644511149
transform 1 0 53452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_581
timestamp 1644511149
transform 1 0 54556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_593
timestamp 1644511149
transform 1 0 55660 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_598
timestamp 1644511149
transform 1 0 56120 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_610
timestamp 1644511149
transform 1 0 57224 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1644511149
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_185
timestamp 1644511149
transform 1 0 18124 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_213
timestamp 1644511149
transform 1 0 20700 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_220
timestamp 1644511149
transform 1 0 21344 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_240
timestamp 1644511149
transform 1 0 23184 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_244
timestamp 1644511149
transform 1 0 23552 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1644511149
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_269
timestamp 1644511149
transform 1 0 25852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_284
timestamp 1644511149
transform 1 0 27232 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_304
timestamp 1644511149
transform 1 0 29072 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_341
timestamp 1644511149
transform 1 0 32476 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_347
timestamp 1644511149
transform 1 0 33028 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_356
timestamp 1644511149
transform 1 0 33856 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_368
timestamp 1644511149
transform 1 0 34960 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_376
timestamp 1644511149
transform 1 0 35696 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_383
timestamp 1644511149
transform 1 0 36340 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_395
timestamp 1644511149
transform 1 0 37444 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_403
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_414
timestamp 1644511149
transform 1 0 39192 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_429
timestamp 1644511149
transform 1 0 40572 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_437
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_445
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_454
timestamp 1644511149
transform 1 0 42872 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_466
timestamp 1644511149
transform 1 0 43976 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_471
timestamp 1644511149
transform 1 0 44436 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_480
timestamp 1644511149
transform 1 0 45264 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_499
timestamp 1644511149
transform 1 0 47012 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_510
timestamp 1644511149
transform 1 0 48024 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_522
timestamp 1644511149
transform 1 0 49128 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_530
timestamp 1644511149
transform 1 0 49864 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_533
timestamp 1644511149
transform 1 0 50140 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_539
timestamp 1644511149
transform 1 0 50692 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_546
timestamp 1644511149
transform 1 0 51336 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_558
timestamp 1644511149
transform 1 0 52440 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_570
timestamp 1644511149
transform 1 0 53544 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_582
timestamp 1644511149
transform 1 0 54648 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_589
timestamp 1644511149
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_601
timestamp 1644511149
transform 1 0 56396 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_610
timestamp 1644511149
transform 1 0 57224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_617
timestamp 1644511149
transform 1 0 57868 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_211
timestamp 1644511149
transform 1 0 20516 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_233
timestamp 1644511149
transform 1 0 22540 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_241
timestamp 1644511149
transform 1 0 23276 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_250
timestamp 1644511149
transform 1 0 24104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_254
timestamp 1644511149
transform 1 0 24472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_260
timestamp 1644511149
transform 1 0 25024 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_264
timestamp 1644511149
transform 1 0 25392 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_268
timestamp 1644511149
transform 1 0 25760 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_285
timestamp 1644511149
transform 1 0 27324 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_290
timestamp 1644511149
transform 1 0 27784 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_310
timestamp 1644511149
transform 1 0 29624 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_330
timestamp 1644511149
transform 1 0 31464 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_345
timestamp 1644511149
transform 1 0 32844 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_357
timestamp 1644511149
transform 1 0 33948 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_369
timestamp 1644511149
transform 1 0 35052 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_387
timestamp 1644511149
transform 1 0 36708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_399
timestamp 1644511149
transform 1 0 37812 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_403
timestamp 1644511149
transform 1 0 38180 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_411
timestamp 1644511149
transform 1 0 38916 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_417
timestamp 1644511149
transform 1 0 39468 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_429
timestamp 1644511149
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_453
timestamp 1644511149
transform 1 0 42780 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_81_468
timestamp 1644511149
transform 1 0 44160 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_479
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_486
timestamp 1644511149
transform 1 0 45816 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_494
timestamp 1644511149
transform 1 0 46552 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_515
timestamp 1644511149
transform 1 0 48484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_527
timestamp 1644511149
transform 1 0 49588 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_533
timestamp 1644511149
transform 1 0 50140 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_544
timestamp 1644511149
transform 1 0 51152 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_556
timestamp 1644511149
transform 1 0 52256 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_561
timestamp 1644511149
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_573
timestamp 1644511149
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_585
timestamp 1644511149
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_597
timestamp 1644511149
transform 1 0 56028 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_605
timestamp 1644511149
transform 1 0 56764 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1644511149
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1644511149
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_620
timestamp 1644511149
transform 1 0 58144 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_624
timestamp 1644511149
transform 1 0 58512 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1644511149
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_177
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_214
timestamp 1644511149
transform 1 0 20792 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_223
timestamp 1644511149
transform 1 0 21620 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_231
timestamp 1644511149
transform 1 0 22356 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_269
timestamp 1644511149
transform 1 0 25852 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_304
timestamp 1644511149
transform 1 0 29072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_316
timestamp 1644511149
transform 1 0 30176 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_326
timestamp 1644511149
transform 1 0 31096 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_353
timestamp 1644511149
transform 1 0 33580 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_372
timestamp 1644511149
transform 1 0 35328 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_380
timestamp 1644511149
transform 1 0 36064 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_385
timestamp 1644511149
transform 1 0 36524 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_397
timestamp 1644511149
transform 1 0 37628 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_409
timestamp 1644511149
transform 1 0 38732 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1644511149
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_428
timestamp 1644511149
transform 1 0 40480 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_436
timestamp 1644511149
transform 1 0 41216 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_442
timestamp 1644511149
transform 1 0 41768 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_451
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_459
timestamp 1644511149
transform 1 0 43332 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_484
timestamp 1644511149
transform 1 0 45632 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_492
timestamp 1644511149
transform 1 0 46368 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_502
timestamp 1644511149
transform 1 0 47288 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_513
timestamp 1644511149
transform 1 0 48300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_524
timestamp 1644511149
transform 1 0 49312 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_539
timestamp 1644511149
transform 1 0 50692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_551
timestamp 1644511149
transform 1 0 51796 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_563
timestamp 1644511149
transform 1 0 52900 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_575
timestamp 1644511149
transform 1 0 54004 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1644511149
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_589
timestamp 1644511149
transform 1 0 55292 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_597
timestamp 1644511149
transform 1 0 56028 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_621
timestamp 1644511149
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1644511149
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1644511149
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1644511149
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1644511149
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1644511149
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1644511149
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1644511149
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_125
timestamp 1644511149
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_137
timestamp 1644511149
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_149
timestamp 1644511149
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1644511149
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1644511149
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_181
timestamp 1644511149
transform 1 0 17756 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_189
timestamp 1644511149
transform 1 0 18492 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_208
timestamp 1644511149
transform 1 0 20240 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_215
timestamp 1644511149
transform 1 0 20884 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1644511149
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_237
timestamp 1644511149
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_257
timestamp 1644511149
transform 1 0 24748 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_265
timestamp 1644511149
transform 1 0 25484 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_272
timestamp 1644511149
transform 1 0 26128 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_289
timestamp 1644511149
transform 1 0 27692 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_293
timestamp 1644511149
transform 1 0 28060 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_306
timestamp 1644511149
transform 1 0 29256 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_314
timestamp 1644511149
transform 1 0 29992 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_321
timestamp 1644511149
transform 1 0 30636 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_325
timestamp 1644511149
transform 1 0 31004 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1644511149
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1644511149
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_343
timestamp 1644511149
transform 1 0 32660 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_355
timestamp 1644511149
transform 1 0 33764 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_375
timestamp 1644511149
transform 1 0 35604 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_387
timestamp 1644511149
transform 1 0 36708 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1644511149
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_400
timestamp 1644511149
transform 1 0 37904 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_412
timestamp 1644511149
transform 1 0 39008 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_424
timestamp 1644511149
transform 1 0 40112 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_432
timestamp 1644511149
transform 1 0 40848 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_436
timestamp 1644511149
transform 1 0 41216 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_442
timestamp 1644511149
transform 1 0 41768 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_449
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_461
timestamp 1644511149
transform 1 0 43516 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_467
timestamp 1644511149
transform 1 0 44068 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_473
timestamp 1644511149
transform 1 0 44620 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_485
timestamp 1644511149
transform 1 0 45724 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_495
timestamp 1644511149
transform 1 0 46644 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1644511149
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_513
timestamp 1644511149
transform 1 0 48300 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_524
timestamp 1644511149
transform 1 0 49312 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_536
timestamp 1644511149
transform 1 0 50416 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_548
timestamp 1644511149
transform 1 0 51520 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_561
timestamp 1644511149
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_573
timestamp 1644511149
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_585
timestamp 1644511149
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_597
timestamp 1644511149
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1644511149
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1644511149
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1644511149
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1644511149
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1644511149
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1644511149
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1644511149
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_97
timestamp 1644511149
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_109
timestamp 1644511149
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_121
timestamp 1644511149
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1644511149
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1644511149
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_153
timestamp 1644511149
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_165
timestamp 1644511149
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_177
timestamp 1644511149
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1644511149
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1644511149
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_197
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_206
timestamp 1644511149
transform 1 0 20056 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_218
timestamp 1644511149
transform 1 0 21160 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_230
timestamp 1644511149
transform 1 0 22264 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_242
timestamp 1644511149
transform 1 0 23368 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_248
timestamp 1644511149
transform 1 0 23920 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_258
timestamp 1644511149
transform 1 0 24840 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_262
timestamp 1644511149
transform 1 0 25208 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_273
timestamp 1644511149
transform 1 0 26220 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_285
timestamp 1644511149
transform 1 0 27324 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_289
timestamp 1644511149
transform 1 0 27692 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_300
timestamp 1644511149
transform 1 0 28704 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_309
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_321
timestamp 1644511149
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_333
timestamp 1644511149
transform 1 0 31740 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_340
timestamp 1644511149
transform 1 0 32384 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_360
timestamp 1644511149
transform 1 0 34224 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_377
timestamp 1644511149
transform 1 0 35788 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_385
timestamp 1644511149
transform 1 0 36524 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_394
timestamp 1644511149
transform 1 0 37352 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_405
timestamp 1644511149
transform 1 0 38364 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_417
timestamp 1644511149
transform 1 0 39468 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_425
timestamp 1644511149
transform 1 0 40204 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_437
timestamp 1644511149
transform 1 0 41308 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_453
timestamp 1644511149
transform 1 0 42780 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_465
timestamp 1644511149
transform 1 0 43884 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_470
timestamp 1644511149
transform 1 0 44344 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_484
timestamp 1644511149
transform 1 0 45632 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_492
timestamp 1644511149
transform 1 0 46368 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_496
timestamp 1644511149
transform 1 0 46736 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_504
timestamp 1644511149
transform 1 0 47472 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_508
timestamp 1644511149
transform 1 0 47840 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_512
timestamp 1644511149
transform 1 0 48208 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_524
timestamp 1644511149
transform 1 0 49312 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_533
timestamp 1644511149
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_545
timestamp 1644511149
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_557
timestamp 1644511149
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_569
timestamp 1644511149
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1644511149
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1644511149
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_589
timestamp 1644511149
transform 1 0 55292 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_597
timestamp 1644511149
transform 1 0 56028 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_621
timestamp 1644511149
transform 1 0 58236 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1644511149
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1644511149
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1644511149
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1644511149
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1644511149
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_76
timestamp 1644511149
transform 1 0 8096 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_101
timestamp 1644511149
transform 1 0 10396 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_109
timestamp 1644511149
transform 1 0 11132 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_113
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_125
timestamp 1644511149
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_137
timestamp 1644511149
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_149
timestamp 1644511149
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1644511149
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1644511149
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_169
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_181
timestamp 1644511149
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_193
timestamp 1644511149
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_205
timestamp 1644511149
transform 1 0 19964 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_85_213
timestamp 1644511149
transform 1 0 20700 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_221
timestamp 1644511149
transform 1 0 21436 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_244
timestamp 1644511149
transform 1 0 23552 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_248
timestamp 1644511149
transform 1 0 23920 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_255
timestamp 1644511149
transform 1 0 24564 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_259
timestamp 1644511149
transform 1 0 24932 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_276
timestamp 1644511149
transform 1 0 26496 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_284
timestamp 1644511149
transform 1 0 27232 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_293
timestamp 1644511149
transform 1 0 28060 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_302
timestamp 1644511149
transform 1 0 28888 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_311
timestamp 1644511149
transform 1 0 29716 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_323
timestamp 1644511149
transform 1 0 30820 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1644511149
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_337
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_349
timestamp 1644511149
transform 1 0 33212 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_353
timestamp 1644511149
transform 1 0 33580 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_361
timestamp 1644511149
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_373
timestamp 1644511149
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1644511149
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1644511149
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_393
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_410
timestamp 1644511149
transform 1 0 38824 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_423
timestamp 1644511149
transform 1 0 40020 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_437
timestamp 1644511149
transform 1 0 41308 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_444
timestamp 1644511149
transform 1 0 41952 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_458
timestamp 1644511149
transform 1 0 43240 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_467
timestamp 1644511149
transform 1 0 44068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_473
timestamp 1644511149
transform 1 0 44620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_481
timestamp 1644511149
transform 1 0 45356 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_493
timestamp 1644511149
transform 1 0 46460 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_501
timestamp 1644511149
transform 1 0 47196 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_85_514
timestamp 1644511149
transform 1 0 48392 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_526
timestamp 1644511149
transform 1 0 49496 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_538
timestamp 1644511149
transform 1 0 50600 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_550
timestamp 1644511149
transform 1 0 51704 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_558
timestamp 1644511149
transform 1 0 52440 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_561
timestamp 1644511149
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_573
timestamp 1644511149
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_585
timestamp 1644511149
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_597
timestamp 1644511149
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1644511149
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1644511149
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1644511149
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1644511149
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1644511149
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1644511149
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_97
timestamp 1644511149
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_109
timestamp 1644511149
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1644511149
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1644511149
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_153
timestamp 1644511149
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_165
timestamp 1644511149
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_177
timestamp 1644511149
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1644511149
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1644511149
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_213
timestamp 1644511149
transform 1 0 20700 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_221
timestamp 1644511149
transform 1 0 21436 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_239
timestamp 1644511149
transform 1 0 23092 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_248
timestamp 1644511149
transform 1 0 23920 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_269
timestamp 1644511149
transform 1 0 25852 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_278
timestamp 1644511149
transform 1 0 26680 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_286
timestamp 1644511149
transform 1 0 27416 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1644511149
transform 1 0 29072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_315
timestamp 1644511149
transform 1 0 30084 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_323
timestamp 1644511149
transform 1 0 30820 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_335
timestamp 1644511149
transform 1 0 31924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_347
timestamp 1644511149
transform 1 0 33028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_359
timestamp 1644511149
transform 1 0 34132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1644511149
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_381
timestamp 1644511149
transform 1 0 36156 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_393
timestamp 1644511149
transform 1 0 37260 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_410
timestamp 1644511149
transform 1 0 38824 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_418
timestamp 1644511149
transform 1 0 39560 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_431
timestamp 1644511149
transform 1 0 40756 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_441
timestamp 1644511149
transform 1 0 41676 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_450
timestamp 1644511149
transform 1 0 42504 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_459
timestamp 1644511149
transform 1 0 43332 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_471
timestamp 1644511149
transform 1 0 44436 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1644511149
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_477
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_489
timestamp 1644511149
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_501
timestamp 1644511149
transform 1 0 47196 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_528
timestamp 1644511149
transform 1 0 49680 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_533
timestamp 1644511149
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_545
timestamp 1644511149
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_557
timestamp 1644511149
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_569
timestamp 1644511149
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1644511149
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1644511149
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_589
timestamp 1644511149
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_601
timestamp 1644511149
transform 1 0 56396 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_607
timestamp 1644511149
transform 1 0 56948 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_611
timestamp 1644511149
transform 1 0 57316 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_618
timestamp 1644511149
transform 1 0 57960 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_624
timestamp 1644511149
transform 1 0 58512 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1644511149
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1644511149
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1644511149
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1644511149
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1644511149
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1644511149
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1644511149
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_113
timestamp 1644511149
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_125
timestamp 1644511149
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_137
timestamp 1644511149
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_149
timestamp 1644511149
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1644511149
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1644511149
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_169
timestamp 1644511149
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_181
timestamp 1644511149
transform 1 0 17756 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_189
timestamp 1644511149
transform 1 0 18492 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_195
timestamp 1644511149
transform 1 0 19044 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_204
timestamp 1644511149
transform 1 0 19872 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_215
timestamp 1644511149
transform 1 0 20884 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1644511149
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_225
timestamp 1644511149
transform 1 0 21804 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_231
timestamp 1644511149
transform 1 0 22356 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_235
timestamp 1644511149
transform 1 0 22724 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_246
timestamp 1644511149
transform 1 0 23736 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_257
timestamp 1644511149
transform 1 0 24748 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_263
timestamp 1644511149
transform 1 0 25300 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_274
timestamp 1644511149
transform 1 0 26312 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_281
timestamp 1644511149
transform 1 0 26956 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_289
timestamp 1644511149
transform 1 0 27692 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_311
timestamp 1644511149
transform 1 0 29716 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_320
timestamp 1644511149
transform 1 0 30544 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_327
timestamp 1644511149
transform 1 0 31188 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1644511149
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_344
timestamp 1644511149
transform 1 0 32752 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_351
timestamp 1644511149
transform 1 0 33396 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_363
timestamp 1644511149
transform 1 0 34500 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_375
timestamp 1644511149
transform 1 0 35604 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_387
timestamp 1644511149
transform 1 0 36708 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1644511149
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_87_393
timestamp 1644511149
transform 1 0 37260 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_412
timestamp 1644511149
transform 1 0 39008 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_420
timestamp 1644511149
transform 1 0 39744 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_429
timestamp 1644511149
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1644511149
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1644511149
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_449
timestamp 1644511149
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_461
timestamp 1644511149
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_473
timestamp 1644511149
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_485
timestamp 1644511149
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1644511149
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1644511149
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_505
timestamp 1644511149
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_517
timestamp 1644511149
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_529
timestamp 1644511149
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_541
timestamp 1644511149
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1644511149
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1644511149
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_561
timestamp 1644511149
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_573
timestamp 1644511149
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_585
timestamp 1644511149
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_597
timestamp 1644511149
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1644511149
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1644511149
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1644511149
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1644511149
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1644511149
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_97
timestamp 1644511149
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_109
timestamp 1644511149
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_121
timestamp 1644511149
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1644511149
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1644511149
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_141
timestamp 1644511149
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_153
timestamp 1644511149
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_165
timestamp 1644511149
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_177
timestamp 1644511149
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_192
timestamp 1644511149
transform 1 0 18768 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_213
timestamp 1644511149
transform 1 0 20700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_225
timestamp 1644511149
transform 1 0 21804 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_232
timestamp 1644511149
transform 1 0 22448 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_244
timestamp 1644511149
transform 1 0 23552 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_88_253
timestamp 1644511149
transform 1 0 24380 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_257
timestamp 1644511149
transform 1 0 24748 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_262
timestamp 1644511149
transform 1 0 25208 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_268
timestamp 1644511149
transform 1 0 25760 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_279
timestamp 1644511149
transform 1 0 26772 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_287
timestamp 1644511149
transform 1 0 27508 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_304
timestamp 1644511149
transform 1 0 29072 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_317
timestamp 1644511149
transform 1 0 30268 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_328
timestamp 1644511149
transform 1 0 31280 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_336
timestamp 1644511149
transform 1 0 32016 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_353
timestamp 1644511149
transform 1 0 33580 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_361
timestamp 1644511149
transform 1 0 34316 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_365
timestamp 1644511149
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_377
timestamp 1644511149
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_389
timestamp 1644511149
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_401
timestamp 1644511149
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1644511149
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1644511149
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_421
timestamp 1644511149
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_433
timestamp 1644511149
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_445
timestamp 1644511149
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_457
timestamp 1644511149
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1644511149
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1644511149
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_477
timestamp 1644511149
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_489
timestamp 1644511149
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_501
timestamp 1644511149
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_513
timestamp 1644511149
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1644511149
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1644511149
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_533
timestamp 1644511149
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_545
timestamp 1644511149
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_557
timestamp 1644511149
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_569
timestamp 1644511149
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1644511149
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1644511149
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_589
timestamp 1644511149
transform 1 0 55292 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_597
timestamp 1644511149
transform 1 0 56028 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_621
timestamp 1644511149
transform 1 0 58236 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1644511149
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1644511149
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1644511149
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1644511149
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1644511149
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1644511149
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1644511149
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1644511149
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_113
timestamp 1644511149
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_125
timestamp 1644511149
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_137
timestamp 1644511149
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_149
timestamp 1644511149
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1644511149
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1644511149
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_169
timestamp 1644511149
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_181
timestamp 1644511149
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_193
timestamp 1644511149
transform 1 0 18860 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_201
timestamp 1644511149
transform 1 0 19596 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_207
timestamp 1644511149
transform 1 0 20148 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_219
timestamp 1644511149
transform 1 0 21252 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1644511149
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_225
timestamp 1644511149
transform 1 0 21804 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_231
timestamp 1644511149
transform 1 0 22356 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_237
timestamp 1644511149
transform 1 0 22908 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_244
timestamp 1644511149
transform 1 0 23552 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_256
timestamp 1644511149
transform 1 0 24656 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_260
timestamp 1644511149
transform 1 0 25024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_274
timestamp 1644511149
transform 1 0 26312 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_281
timestamp 1644511149
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_293
timestamp 1644511149
transform 1 0 28060 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_297
timestamp 1644511149
transform 1 0 28428 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_314
timestamp 1644511149
transform 1 0 29992 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_323
timestamp 1644511149
transform 1 0 30820 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_332
timestamp 1644511149
transform 1 0 31648 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_353
timestamp 1644511149
transform 1 0 33580 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_363
timestamp 1644511149
transform 1 0 34500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_375
timestamp 1644511149
transform 1 0 35604 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_387
timestamp 1644511149
transform 1 0 36708 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1644511149
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_393
timestamp 1644511149
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_405
timestamp 1644511149
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_417
timestamp 1644511149
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_429
timestamp 1644511149
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1644511149
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1644511149
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_449
timestamp 1644511149
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_461
timestamp 1644511149
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_473
timestamp 1644511149
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_485
timestamp 1644511149
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1644511149
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1644511149
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_505
timestamp 1644511149
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_517
timestamp 1644511149
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_529
timestamp 1644511149
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_541
timestamp 1644511149
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1644511149
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1644511149
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_561
timestamp 1644511149
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_573
timestamp 1644511149
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_585
timestamp 1644511149
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_597
timestamp 1644511149
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1644511149
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1644511149
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1644511149
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1644511149
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1644511149
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_97
timestamp 1644511149
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_109
timestamp 1644511149
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_121
timestamp 1644511149
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1644511149
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1644511149
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_141
timestamp 1644511149
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_153
timestamp 1644511149
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_165
timestamp 1644511149
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_177
timestamp 1644511149
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1644511149
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1644511149
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_213
timestamp 1644511149
transform 1 0 20700 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_221
timestamp 1644511149
transform 1 0 21436 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_226
timestamp 1644511149
transform 1 0 21896 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_235
timestamp 1644511149
transform 1 0 22724 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1644511149
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1644511149
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_253
timestamp 1644511149
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_265
timestamp 1644511149
transform 1 0 25484 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_271
timestamp 1644511149
transform 1 0 26036 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_283
timestamp 1644511149
transform 1 0 27140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_295
timestamp 1644511149
transform 1 0 28244 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_304
timestamp 1644511149
transform 1 0 29072 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_309
timestamp 1644511149
transform 1 0 29532 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_316
timestamp 1644511149
transform 1 0 30176 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_323
timestamp 1644511149
transform 1 0 30820 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_332
timestamp 1644511149
transform 1 0 31648 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_352
timestamp 1644511149
transform 1 0 33488 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_359
timestamp 1644511149
transform 1 0 34132 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1644511149
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_365
timestamp 1644511149
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_377
timestamp 1644511149
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_389
timestamp 1644511149
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_401
timestamp 1644511149
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1644511149
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1644511149
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_421
timestamp 1644511149
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_433
timestamp 1644511149
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_445
timestamp 1644511149
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_457
timestamp 1644511149
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1644511149
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1644511149
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_477
timestamp 1644511149
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_489
timestamp 1644511149
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_501
timestamp 1644511149
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_513
timestamp 1644511149
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1644511149
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1644511149
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_533
timestamp 1644511149
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_545
timestamp 1644511149
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_557
timestamp 1644511149
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_569
timestamp 1644511149
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1644511149
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1644511149
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_589
timestamp 1644511149
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_601
timestamp 1644511149
transform 1 0 56396 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_610
timestamp 1644511149
transform 1 0 57224 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_617
timestamp 1644511149
transform 1 0 57868 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_91_3
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_11
timestamp 1644511149
transform 1 0 2116 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_33
timestamp 1644511149
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1644511149
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1644511149
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1644511149
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1644511149
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_113
timestamp 1644511149
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_125
timestamp 1644511149
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_137
timestamp 1644511149
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_149
timestamp 1644511149
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1644511149
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1644511149
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_169
timestamp 1644511149
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_181
timestamp 1644511149
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_193
timestamp 1644511149
transform 1 0 18860 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_200
timestamp 1644511149
transform 1 0 19504 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_209
timestamp 1644511149
transform 1 0 20332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_221
timestamp 1644511149
transform 1 0 21436 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_91_225
timestamp 1644511149
transform 1 0 21804 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_242
timestamp 1644511149
transform 1 0 23368 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_253
timestamp 1644511149
transform 1 0 24380 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_259
timestamp 1644511149
transform 1 0 24932 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_276
timestamp 1644511149
transform 1 0 26496 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_284
timestamp 1644511149
transform 1 0 27232 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_296
timestamp 1644511149
transform 1 0 28336 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_308
timestamp 1644511149
transform 1 0 29440 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_91_332
timestamp 1644511149
transform 1 0 31648 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_342
timestamp 1644511149
transform 1 0 32568 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_349
timestamp 1644511149
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_361
timestamp 1644511149
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_373
timestamp 1644511149
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1644511149
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1644511149
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_393
timestamp 1644511149
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_405
timestamp 1644511149
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_417
timestamp 1644511149
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_429
timestamp 1644511149
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1644511149
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1644511149
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_449
timestamp 1644511149
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_461
timestamp 1644511149
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_473
timestamp 1644511149
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_485
timestamp 1644511149
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1644511149
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1644511149
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_505
timestamp 1644511149
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_517
timestamp 1644511149
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_529
timestamp 1644511149
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_541
timestamp 1644511149
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1644511149
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1644511149
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_561
timestamp 1644511149
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_573
timestamp 1644511149
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_585
timestamp 1644511149
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_597
timestamp 1644511149
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1644511149
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1644511149
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1644511149
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_92_3
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_11
timestamp 1644511149
transform 1 0 2116 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_16
timestamp 1644511149
transform 1 0 2576 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_23
timestamp 1644511149
transform 1 0 3220 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1644511149
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_32
timestamp 1644511149
transform 1 0 4048 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_44
timestamp 1644511149
transform 1 0 5152 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_56
timestamp 1644511149
transform 1 0 6256 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_68
timestamp 1644511149
transform 1 0 7360 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_80
timestamp 1644511149
transform 1 0 8464 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_97
timestamp 1644511149
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_109
timestamp 1644511149
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_121
timestamp 1644511149
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1644511149
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1644511149
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_141
timestamp 1644511149
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_153
timestamp 1644511149
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_165
timestamp 1644511149
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_177
timestamp 1644511149
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1644511149
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1644511149
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_197
timestamp 1644511149
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_209
timestamp 1644511149
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_224
timestamp 1644511149
transform 1 0 21712 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_244
timestamp 1644511149
transform 1 0 23552 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_253
timestamp 1644511149
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_281
timestamp 1644511149
transform 1 0 26956 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_293
timestamp 1644511149
transform 1 0 28060 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_305
timestamp 1644511149
transform 1 0 29164 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_309
timestamp 1644511149
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_321
timestamp 1644511149
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_333
timestamp 1644511149
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_345
timestamp 1644511149
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1644511149
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1644511149
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_365
timestamp 1644511149
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_377
timestamp 1644511149
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_389
timestamp 1644511149
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_401
timestamp 1644511149
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1644511149
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1644511149
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_421
timestamp 1644511149
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_433
timestamp 1644511149
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_445
timestamp 1644511149
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_457
timestamp 1644511149
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1644511149
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1644511149
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_477
timestamp 1644511149
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_489
timestamp 1644511149
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_501
timestamp 1644511149
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_513
timestamp 1644511149
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1644511149
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1644511149
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_533
timestamp 1644511149
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_545
timestamp 1644511149
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_557
timestamp 1644511149
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_569
timestamp 1644511149
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1644511149
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1644511149
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_589
timestamp 1644511149
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_601
timestamp 1644511149
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_613
timestamp 1644511149
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_3
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_30
timestamp 1644511149
transform 1 0 3864 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_42
timestamp 1644511149
transform 1 0 4968 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1644511149
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_93
timestamp 1644511149
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1644511149
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1644511149
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_113
timestamp 1644511149
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_125
timestamp 1644511149
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_137
timestamp 1644511149
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_149
timestamp 1644511149
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1644511149
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1644511149
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_169
timestamp 1644511149
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_181
timestamp 1644511149
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_193
timestamp 1644511149
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_205
timestamp 1644511149
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1644511149
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1644511149
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_241
timestamp 1644511149
transform 1 0 23276 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_250
timestamp 1644511149
transform 1 0 24104 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_262
timestamp 1644511149
transform 1 0 25208 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_267
timestamp 1644511149
transform 1 0 25668 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_276
timestamp 1644511149
transform 1 0 26496 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_287
timestamp 1644511149
transform 1 0 27508 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_294
timestamp 1644511149
transform 1 0 28152 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_306
timestamp 1644511149
transform 1 0 29256 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_318
timestamp 1644511149
transform 1 0 30360 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_330
timestamp 1644511149
transform 1 0 31464 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_337
timestamp 1644511149
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_349
timestamp 1644511149
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_361
timestamp 1644511149
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_373
timestamp 1644511149
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1644511149
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1644511149
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_393
timestamp 1644511149
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_405
timestamp 1644511149
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_417
timestamp 1644511149
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_429
timestamp 1644511149
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1644511149
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1644511149
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_449
timestamp 1644511149
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_461
timestamp 1644511149
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_473
timestamp 1644511149
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_485
timestamp 1644511149
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1644511149
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1644511149
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_505
timestamp 1644511149
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_517
timestamp 1644511149
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_529
timestamp 1644511149
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_541
timestamp 1644511149
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1644511149
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1644511149
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_561
timestamp 1644511149
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_573
timestamp 1644511149
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_585
timestamp 1644511149
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_597
timestamp 1644511149
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1644511149
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1644511149
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_620
timestamp 1644511149
transform 1 0 58144 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_624
timestamp 1644511149
transform 1 0 58512 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1644511149
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_13
timestamp 1644511149
transform 1 0 2300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_25
timestamp 1644511149
transform 1 0 3404 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1644511149
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1644511149
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1644511149
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_97
timestamp 1644511149
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_109
timestamp 1644511149
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_121
timestamp 1644511149
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1644511149
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1644511149
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_141
timestamp 1644511149
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_153
timestamp 1644511149
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_165
timestamp 1644511149
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_177
timestamp 1644511149
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1644511149
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1644511149
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_197
timestamp 1644511149
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_209
timestamp 1644511149
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_221
timestamp 1644511149
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_238
timestamp 1644511149
transform 1 0 23000 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1644511149
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_253
timestamp 1644511149
transform 1 0 24380 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_94_277
timestamp 1644511149
transform 1 0 26588 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_288
timestamp 1644511149
transform 1 0 27600 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_94_304
timestamp 1644511149
transform 1 0 29072 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_325
timestamp 1644511149
transform 1 0 31004 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_337
timestamp 1644511149
transform 1 0 32108 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_349
timestamp 1644511149
transform 1 0 33212 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_361
timestamp 1644511149
transform 1 0 34316 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_365
timestamp 1644511149
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_377
timestamp 1644511149
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_389
timestamp 1644511149
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_401
timestamp 1644511149
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1644511149
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1644511149
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_421
timestamp 1644511149
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_433
timestamp 1644511149
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_445
timestamp 1644511149
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_457
timestamp 1644511149
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1644511149
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1644511149
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_477
timestamp 1644511149
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_489
timestamp 1644511149
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_501
timestamp 1644511149
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_513
timestamp 1644511149
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1644511149
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1644511149
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_533
timestamp 1644511149
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_545
timestamp 1644511149
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_557
timestamp 1644511149
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_569
timestamp 1644511149
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1644511149
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1644511149
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_589
timestamp 1644511149
transform 1 0 55292 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_597
timestamp 1644511149
transform 1 0 56028 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_621
timestamp 1644511149
transform 1 0 58236 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1644511149
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1644511149
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_39
timestamp 1644511149
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1644511149
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1644511149
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1644511149
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1644511149
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_93
timestamp 1644511149
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1644511149
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1644511149
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_113
timestamp 1644511149
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_125
timestamp 1644511149
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_137
timestamp 1644511149
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_149
timestamp 1644511149
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1644511149
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1644511149
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_169
timestamp 1644511149
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_181
timestamp 1644511149
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_193
timestamp 1644511149
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_205
timestamp 1644511149
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1644511149
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1644511149
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_225
timestamp 1644511149
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_237
timestamp 1644511149
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_249
timestamp 1644511149
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_261
timestamp 1644511149
transform 1 0 25116 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_95_274
timestamp 1644511149
transform 1 0 26312 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_95_281
timestamp 1644511149
transform 1 0 26956 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_289
timestamp 1644511149
transform 1 0 27692 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_295
timestamp 1644511149
transform 1 0 28244 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_306
timestamp 1644511149
transform 1 0 29256 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_313
timestamp 1644511149
transform 1 0 29900 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_325
timestamp 1644511149
transform 1 0 31004 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_333
timestamp 1644511149
transform 1 0 31740 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_337
timestamp 1644511149
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_349
timestamp 1644511149
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_361
timestamp 1644511149
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_373
timestamp 1644511149
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1644511149
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1644511149
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_393
timestamp 1644511149
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_405
timestamp 1644511149
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_417
timestamp 1644511149
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_429
timestamp 1644511149
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1644511149
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1644511149
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_449
timestamp 1644511149
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_461
timestamp 1644511149
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_473
timestamp 1644511149
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_485
timestamp 1644511149
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1644511149
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1644511149
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_505
timestamp 1644511149
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_517
timestamp 1644511149
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_529
timestamp 1644511149
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_541
timestamp 1644511149
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1644511149
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1644511149
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_561
timestamp 1644511149
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_573
timestamp 1644511149
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_585
timestamp 1644511149
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_597
timestamp 1644511149
transform 1 0 56028 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_602
timestamp 1644511149
transform 1 0 56488 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1644511149
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1644511149
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_620
timestamp 1644511149
transform 1 0 58144 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_624
timestamp 1644511149
transform 1 0 58512 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1644511149
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_18
timestamp 1644511149
transform 1 0 2760 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_26
timestamp 1644511149
transform 1 0 3496 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_32
timestamp 1644511149
transform 1 0 4048 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_44
timestamp 1644511149
transform 1 0 5152 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_56
timestamp 1644511149
transform 1 0 6256 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_68
timestamp 1644511149
transform 1 0 7360 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_80
timestamp 1644511149
transform 1 0 8464 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_97
timestamp 1644511149
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_109
timestamp 1644511149
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_121
timestamp 1644511149
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1644511149
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1644511149
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_141
timestamp 1644511149
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_153
timestamp 1644511149
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_165
timestamp 1644511149
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_177
timestamp 1644511149
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1644511149
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1644511149
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_200
timestamp 1644511149
transform 1 0 19504 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_96_222
timestamp 1644511149
transform 1 0 21528 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_234
timestamp 1644511149
transform 1 0 22632 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_246
timestamp 1644511149
transform 1 0 23736 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_96_253
timestamp 1644511149
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_265
timestamp 1644511149
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_277
timestamp 1644511149
transform 1 0 26588 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_283
timestamp 1644511149
transform 1 0 27140 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_289
timestamp 1644511149
transform 1 0 27692 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_299
timestamp 1644511149
transform 1 0 28612 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1644511149
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_325
timestamp 1644511149
transform 1 0 31004 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_337
timestamp 1644511149
transform 1 0 32108 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_345
timestamp 1644511149
transform 1 0 32844 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_352
timestamp 1644511149
transform 1 0 33488 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_365
timestamp 1644511149
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_377
timestamp 1644511149
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_389
timestamp 1644511149
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_401
timestamp 1644511149
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1644511149
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1644511149
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_421
timestamp 1644511149
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_433
timestamp 1644511149
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_445
timestamp 1644511149
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_457
timestamp 1644511149
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1644511149
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1644511149
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_477
timestamp 1644511149
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_489
timestamp 1644511149
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_501
timestamp 1644511149
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_513
timestamp 1644511149
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1644511149
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1644511149
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_533
timestamp 1644511149
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_545
timestamp 1644511149
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_557
timestamp 1644511149
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_569
timestamp 1644511149
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1644511149
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1644511149
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_589
timestamp 1644511149
transform 1 0 55292 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_597
timestamp 1644511149
transform 1 0 56028 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_621
timestamp 1644511149
transform 1 0 58236 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_3
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_11
timestamp 1644511149
transform 1 0 2116 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_34
timestamp 1644511149
transform 1 0 4232 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_46
timestamp 1644511149
transform 1 0 5336 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_54
timestamp 1644511149
transform 1 0 6072 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_93
timestamp 1644511149
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1644511149
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1644511149
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_113
timestamp 1644511149
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_125
timestamp 1644511149
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_137
timestamp 1644511149
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_149
timestamp 1644511149
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1644511149
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1644511149
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_169
timestamp 1644511149
transform 1 0 16652 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_177
timestamp 1644511149
transform 1 0 17388 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_201
timestamp 1644511149
transform 1 0 19596 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_213
timestamp 1644511149
transform 1 0 20700 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_220
timestamp 1644511149
transform 1 0 21344 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_241
timestamp 1644511149
transform 1 0 23276 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_253
timestamp 1644511149
transform 1 0 24380 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_261
timestamp 1644511149
transform 1 0 25116 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_267
timestamp 1644511149
transform 1 0 25668 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_276
timestamp 1644511149
transform 1 0 26496 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_281
timestamp 1644511149
transform 1 0 26956 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_285
timestamp 1644511149
transform 1 0 27324 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_302
timestamp 1644511149
transform 1 0 28888 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_309
timestamp 1644511149
transform 1 0 29532 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_321
timestamp 1644511149
transform 1 0 30636 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_333
timestamp 1644511149
transform 1 0 31740 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_337
timestamp 1644511149
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_349
timestamp 1644511149
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_361
timestamp 1644511149
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_373
timestamp 1644511149
transform 1 0 35420 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_97_384
timestamp 1644511149
transform 1 0 36432 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_393
timestamp 1644511149
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_405
timestamp 1644511149
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_417
timestamp 1644511149
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_429
timestamp 1644511149
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1644511149
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1644511149
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_449
timestamp 1644511149
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_461
timestamp 1644511149
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_473
timestamp 1644511149
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_485
timestamp 1644511149
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1644511149
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1644511149
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_505
timestamp 1644511149
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_517
timestamp 1644511149
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_529
timestamp 1644511149
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_541
timestamp 1644511149
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1644511149
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1644511149
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_561
timestamp 1644511149
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_573
timestamp 1644511149
transform 1 0 53820 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_97_584
timestamp 1644511149
transform 1 0 54832 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_590
timestamp 1644511149
transform 1 0 55384 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_612
timestamp 1644511149
transform 1 0 57408 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_620
timestamp 1644511149
transform 1 0 58144 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_624
timestamp 1644511149
transform 1 0 58512 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_12
timestamp 1644511149
transform 1 0 2208 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_19
timestamp 1644511149
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1644511149
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_50
timestamp 1644511149
transform 1 0 5704 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_62
timestamp 1644511149
transform 1 0 6808 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_71
timestamp 1644511149
transform 1 0 7636 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1644511149
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_88
timestamp 1644511149
transform 1 0 9200 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_100
timestamp 1644511149
transform 1 0 10304 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_112
timestamp 1644511149
transform 1 0 11408 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_124
timestamp 1644511149
transform 1 0 12512 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_128
timestamp 1644511149
transform 1 0 12880 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_132
timestamp 1644511149
transform 1 0 13248 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_98_141
timestamp 1644511149
transform 1 0 14076 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_149
timestamp 1644511149
transform 1 0 14812 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_155
timestamp 1644511149
transform 1 0 15364 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_180
timestamp 1644511149
transform 1 0 17664 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_192
timestamp 1644511149
transform 1 0 18768 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_200
timestamp 1644511149
transform 1 0 19504 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_208
timestamp 1644511149
transform 1 0 20240 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_212
timestamp 1644511149
transform 1 0 20608 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_219
timestamp 1644511149
transform 1 0 21252 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_223
timestamp 1644511149
transform 1 0 21620 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_229
timestamp 1644511149
transform 1 0 22172 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_236
timestamp 1644511149
transform 1 0 22816 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_248
timestamp 1644511149
transform 1 0 23920 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_253
timestamp 1644511149
transform 1 0 24380 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_98_275
timestamp 1644511149
transform 1 0 26404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_281
timestamp 1644511149
transform 1 0 26956 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_298
timestamp 1644511149
transform 1 0 28520 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_306
timestamp 1644511149
transform 1 0 29256 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_309
timestamp 1644511149
transform 1 0 29532 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_313
timestamp 1644511149
transform 1 0 29900 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_335
timestamp 1644511149
transform 1 0 31924 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_342
timestamp 1644511149
transform 1 0 32568 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_351
timestamp 1644511149
transform 1 0 33396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1644511149
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_365
timestamp 1644511149
transform 1 0 34684 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_372
timestamp 1644511149
transform 1 0 35328 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_397
timestamp 1644511149
transform 1 0 37628 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_409
timestamp 1644511149
transform 1 0 38732 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_417
timestamp 1644511149
transform 1 0 39468 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_421
timestamp 1644511149
transform 1 0 39836 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_98_426
timestamp 1644511149
transform 1 0 40296 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_438
timestamp 1644511149
transform 1 0 41400 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_446
timestamp 1644511149
transform 1 0 42136 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_98_470
timestamp 1644511149
transform 1 0 44344 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_477
timestamp 1644511149
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_489
timestamp 1644511149
transform 1 0 46092 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_511
timestamp 1644511149
transform 1 0 48116 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_523
timestamp 1644511149
transform 1 0 49220 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1644511149
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_536
timestamp 1644511149
transform 1 0 50416 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_548
timestamp 1644511149
transform 1 0 51520 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_560
timestamp 1644511149
transform 1 0 52624 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_584
timestamp 1644511149
transform 1 0 54832 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_589
timestamp 1644511149
transform 1 0 55292 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_596
timestamp 1644511149
transform 1 0 55936 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_621
timestamp 1644511149
transform 1 0 58236 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_3
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_30
timestamp 1644511149
transform 1 0 3864 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_37
timestamp 1644511149
transform 1 0 4508 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_49
timestamp 1644511149
transform 1 0 5612 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1644511149
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_78
timestamp 1644511149
transform 1 0 8280 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_103
timestamp 1644511149
transform 1 0 10580 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1644511149
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_113
timestamp 1644511149
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_125
timestamp 1644511149
transform 1 0 12604 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_131
timestamp 1644511149
transform 1 0 13156 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_153
timestamp 1644511149
transform 1 0 15180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_165
timestamp 1644511149
transform 1 0 16284 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_99_169
timestamp 1644511149
transform 1 0 16652 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_191
timestamp 1644511149
transform 1 0 18676 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_216
timestamp 1644511149
transform 1 0 20976 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_99_230
timestamp 1644511149
transform 1 0 22264 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_254
timestamp 1644511149
transform 1 0 24472 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_266
timestamp 1644511149
transform 1 0 25576 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_270
timestamp 1644511149
transform 1 0 25944 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_276
timestamp 1644511149
transform 1 0 26496 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_286
timestamp 1644511149
transform 1 0 27416 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_99_313
timestamp 1644511149
transform 1 0 29900 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_321
timestamp 1644511149
transform 1 0 30636 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_326
timestamp 1644511149
transform 1 0 31096 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_334
timestamp 1644511149
transform 1 0 31832 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_358
timestamp 1644511149
transform 1 0 34040 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_370
timestamp 1644511149
transform 1 0 35144 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_376
timestamp 1644511149
transform 1 0 35696 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_380
timestamp 1644511149
transform 1 0 36064 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_393
timestamp 1644511149
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_405
timestamp 1644511149
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_417
timestamp 1644511149
transform 1 0 39468 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_440
timestamp 1644511149
transform 1 0 41584 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_449
timestamp 1644511149
transform 1 0 42412 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_472
timestamp 1644511149
transform 1 0 44528 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_484
timestamp 1644511149
transform 1 0 45632 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_492
timestamp 1644511149
transform 1 0 46368 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_498
timestamp 1644511149
transform 1 0 46920 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_505
timestamp 1644511149
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_517
timestamp 1644511149
transform 1 0 48668 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_525
timestamp 1644511149
transform 1 0 49404 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_547
timestamp 1644511149
transform 1 0 51428 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1644511149
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_561
timestamp 1644511149
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_573
timestamp 1644511149
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_585
timestamp 1644511149
transform 1 0 54924 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_612
timestamp 1644511149
transform 1 0 57408 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_620
timestamp 1644511149
transform 1 0 58144 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_624
timestamp 1644511149
transform 1 0 58512 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_3
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_9
timestamp 1644511149
transform 1 0 1932 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_13
timestamp 1644511149
transform 1 0 2300 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_20
timestamp 1644511149
transform 1 0 2944 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_100_50
timestamp 1644511149
transform 1 0 5704 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_100_59
timestamp 1644511149
transform 1 0 6532 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_67
timestamp 1644511149
transform 1 0 7268 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_72
timestamp 1644511149
transform 1 0 7728 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_97
timestamp 1644511149
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_109
timestamp 1644511149
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_121
timestamp 1644511149
transform 1 0 12236 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_129
timestamp 1644511149
transform 1 0 12972 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_135
timestamp 1644511149
transform 1 0 13524 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1644511149
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_141
timestamp 1644511149
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_153
timestamp 1644511149
transform 1 0 15180 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_159
timestamp 1644511149
transform 1 0 15732 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_163
timestamp 1644511149
transform 1 0 16100 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_175
timestamp 1644511149
transform 1 0 17204 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_180
timestamp 1644511149
transform 1 0 17664 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_187
timestamp 1644511149
transform 1 0 18308 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1644511149
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_197
timestamp 1644511149
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_209
timestamp 1644511149
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_221
timestamp 1644511149
transform 1 0 21436 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_229
timestamp 1644511149
transform 1 0 22172 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_234
timestamp 1644511149
transform 1 0 22632 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_246
timestamp 1644511149
transform 1 0 23736 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_100_253
timestamp 1644511149
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_265
timestamp 1644511149
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_277
timestamp 1644511149
transform 1 0 26588 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_281
timestamp 1644511149
transform 1 0 26956 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_285
timestamp 1644511149
transform 1 0 27324 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_292
timestamp 1644511149
transform 1 0 27968 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_299
timestamp 1644511149
transform 1 0 28612 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1644511149
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_309
timestamp 1644511149
transform 1 0 29532 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_313
timestamp 1644511149
transform 1 0 29900 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_317
timestamp 1644511149
transform 1 0 30268 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_324
timestamp 1644511149
transform 1 0 30912 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_349
timestamp 1644511149
transform 1 0 33212 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_361
timestamp 1644511149
transform 1 0 34316 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_365
timestamp 1644511149
transform 1 0 34684 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_373
timestamp 1644511149
transform 1 0 35420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_396
timestamp 1644511149
transform 1 0 37536 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_408
timestamp 1644511149
transform 1 0 38640 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_424
timestamp 1644511149
transform 1 0 40112 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_436
timestamp 1644511149
transform 1 0 41216 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_444
timestamp 1644511149
transform 1 0 41952 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_448
timestamp 1644511149
transform 1 0 42320 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_455
timestamp 1644511149
transform 1 0 42964 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_467
timestamp 1644511149
transform 1 0 44068 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1644511149
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_477
timestamp 1644511149
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_489
timestamp 1644511149
transform 1 0 46092 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_494
timestamp 1644511149
transform 1 0 46552 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_506
timestamp 1644511149
transform 1 0 47656 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_518
timestamp 1644511149
transform 1 0 48760 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_530
timestamp 1644511149
transform 1 0 49864 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_536
timestamp 1644511149
transform 1 0 50416 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_548
timestamp 1644511149
transform 1 0 51520 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_560
timestamp 1644511149
transform 1 0 52624 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_572
timestamp 1644511149
transform 1 0 53728 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_584
timestamp 1644511149
transform 1 0 54832 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_589
timestamp 1644511149
transform 1 0 55292 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_596
timestamp 1644511149
transform 1 0 55936 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1644511149
transform 1 0 58236 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_13
timestamp 1644511149
transform 1 0 2300 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_20
timestamp 1644511149
transform 1 0 2944 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_29
timestamp 1644511149
transform 1 0 3772 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_33
timestamp 1644511149
transform 1 0 4140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_45
timestamp 1644511149
transform 1 0 5244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1644511149
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_85
timestamp 1644511149
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_97
timestamp 1644511149
transform 1 0 10028 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_104
timestamp 1644511149
transform 1 0 10672 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_113
timestamp 1644511149
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_125
timestamp 1644511149
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 1644511149
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_141
timestamp 1644511149
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_153
timestamp 1644511149
transform 1 0 15180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_165
timestamp 1644511149
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_169
timestamp 1644511149
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_184
timestamp 1644511149
transform 1 0 18032 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_197
timestamp 1644511149
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_209
timestamp 1644511149
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1644511149
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_225
timestamp 1644511149
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_237
timestamp 1644511149
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1644511149
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_253
timestamp 1644511149
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_265
timestamp 1644511149
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1644511149
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_281
timestamp 1644511149
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_293
timestamp 1644511149
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1644511149
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_309
timestamp 1644511149
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_321
timestamp 1644511149
transform 1 0 30636 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_327
timestamp 1644511149
transform 1 0 31188 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_331
timestamp 1644511149
transform 1 0 31556 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1644511149
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_340
timestamp 1644511149
transform 1 0 32384 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_352
timestamp 1644511149
transform 1 0 33488 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_356
timestamp 1644511149
transform 1 0 33856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_101_365
timestamp 1644511149
transform 1 0 34684 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_373
timestamp 1644511149
transform 1 0 35420 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_379
timestamp 1644511149
transform 1 0 35972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1644511149
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_393
timestamp 1644511149
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_405
timestamp 1644511149
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1644511149
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_421
timestamp 1644511149
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_433
timestamp 1644511149
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1644511149
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_449
timestamp 1644511149
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_461
timestamp 1644511149
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1644511149
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_477
timestamp 1644511149
transform 1 0 44988 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_489
timestamp 1644511149
transform 1 0 46092 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_501
timestamp 1644511149
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_505
timestamp 1644511149
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_517
timestamp 1644511149
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1644511149
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_533
timestamp 1644511149
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_545
timestamp 1644511149
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1644511149
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_561
timestamp 1644511149
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_573
timestamp 1644511149
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1644511149
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_589
timestamp 1644511149
transform 1 0 55292 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_598
timestamp 1644511149
transform 1 0 56120 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_605
timestamp 1644511149
transform 1 0 56764 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_612
timestamp 1644511149
transform 1 0 57408 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_620
timestamp 1644511149
transform 1 0 58144 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_624
timestamp 1644511149
transform 1 0 58512 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1644511149
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1644511149
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1644511149
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1644511149
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1644511149
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1644511149
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1644511149
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1644511149
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1644511149
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1644511149
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1644511149
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1644511149
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1644511149
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1644511149
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1644511149
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1644511149
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1644511149
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1644511149
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1644511149
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1644511149
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1644511149
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1644511149
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1644511149
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1644511149
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1644511149
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1644511149
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1644511149
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1644511149
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1644511149
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1644511149
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1644511149
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1644511149
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1644511149
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1644511149
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1644511149
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1644511149
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1644511149
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1644511149
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1644511149
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1644511149
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1644511149
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1644511149
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1644511149
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1644511149
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1644511149
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1644511149
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1644511149
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1644511149
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1644511149
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1644511149
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1644511149
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1644511149
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1644511149
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1644511149
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1644511149
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1644511149
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1644511149
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1644511149
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1644511149
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1644511149
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1644511149
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1644511149
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1644511149
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1644511149
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1644511149
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1644511149
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1644511149
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1644511149
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1644511149
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1644511149
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1644511149
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1644511149
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1644511149
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1644511149
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1644511149
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1644511149
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1644511149
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1644511149
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1644511149
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1644511149
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1644511149
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1644511149
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1644511149
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1644511149
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1644511149
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1644511149
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1644511149
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1644511149
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1644511149
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1644511149
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1644511149
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1644511149
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1644511149
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1644511149
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1644511149
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1644511149
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1644511149
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1644511149
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1644511149
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1644511149
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1644511149
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1644511149
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1644511149
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1644511149
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1644511149
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1644511149
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1644511149
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1644511149
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1644511149
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1644511149
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1644511149
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1644511149
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1644511149
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1644511149
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1644511149
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1644511149
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1644511149
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1644511149
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1644511149
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1644511149
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1644511149
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1644511149
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1644511149
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1644511149
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1644511149
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1644511149
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1644511149
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1644511149
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1644511149
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1644511149
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1644511149
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1644511149
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1644511149
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1644511149
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1644511149
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1644511149
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1644511149
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1644511149
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1644511149
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1644511149
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1644511149
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1644511149
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1644511149
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1644511149
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1644511149
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1644511149
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1644511149
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1644511149
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1644511149
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1644511149
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1644511149
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1644511149
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1644511149
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1644511149
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1644511149
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1644511149
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1644511149
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1644511149
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1644511149
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1644511149
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1644511149
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1644511149
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _1174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _1175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  _1176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 55568 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1644511149
transform 1 0 56856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1644511149
transform 1 0 55660 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1644511149
transform 1 0 40020 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1182_
timestamp 1644511149
transform 1 0 4232 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1644511149
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1644511149
transform 1 0 56856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1644511149
transform 1 0 28336 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1644511149
transform 1 0 57868 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1188_
timestamp 1644511149
transform 1 0 7636 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8648 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1190_
timestamp 1644511149
transform 1 0 2300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1644511149
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1644511149
transform 1 0 2300 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1194_
timestamp 1644511149
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1196_
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1197_
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198_
timestamp 1644511149
transform 1 0 56856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1199_
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 56856 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  _1201_
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1644511149
transform 1 0 57868 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1644511149
transform 1 0 56856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1644511149
transform 1 0 56856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1644511149
transform 1 0 7360 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1207_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1644511149
transform 1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 1644511149
transform 1 0 46644 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1644511149
transform 1 0 17388 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1644511149
transform 1 0 56304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1212_
timestamp 1644511149
transform 1 0 2576 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1213_
timestamp 1644511149
transform 1 0 8648 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1216_
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1644511149
transform 1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1218_
timestamp 1644511149
transform 1 0 56856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1219_
timestamp 1644511149
transform 1 0 28520 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1644511149
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1222_
timestamp 1644511149
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1223_
timestamp 1644511149
transform 1 0 29532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1644511149
transform 1 0 30360 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1644511149
transform 1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1226_
timestamp 1644511149
transform 1 0 29624 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1227_
timestamp 1644511149
transform 1 0 31096 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1228_
timestamp 1644511149
transform 1 0 7820 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1644511149
transform 1 0 19228 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1231_
timestamp 1644511149
transform 1 0 56212 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1232_
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1233_
timestamp 1644511149
transform 1 0 30820 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1234_
timestamp 1644511149
transform 1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1644511149
transform 1 0 30636 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1236_
timestamp 1644511149
transform 1 0 54832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1237_
timestamp 1644511149
transform 1 0 50140 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1238_
timestamp 1644511149
transform 1 0 30452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1239_
timestamp 1644511149
transform 1 0 56856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1240_
timestamp 1644511149
transform 1 0 31096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1241_
timestamp 1644511149
transform 1 0 35052 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1242_
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1644511149
transform 1 0 49956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1244_
timestamp 1644511149
transform 1 0 29716 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1245_
timestamp 1644511149
transform 1 0 57224 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1246_
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1247_
timestamp 1644511149
transform 1 0 4232 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1248_
timestamp 1644511149
transform 1 0 56948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1249_
timestamp 1644511149
transform 1 0 15088 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _1251_
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1254_
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1256_
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1257_
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1258_
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1259_
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1644511149
transform 1 0 54556 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1261_
timestamp 1644511149
transform 1 0 56580 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1262_
timestamp 1644511149
transform 1 0 57040 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1263_
timestamp 1644511149
transform 1 0 19504 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1264_
timestamp 1644511149
transform 1 0 2392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1644511149
transform 1 0 2392 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1266_
timestamp 1644511149
transform 1 0 57040 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1644511149
transform 1 0 56948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1268_
timestamp 1644511149
transform 1 0 12972 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1269_
timestamp 1644511149
transform 1 0 19412 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1270_
timestamp 1644511149
transform 1 0 57040 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1271_
timestamp 1644511149
transform 1 0 57040 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1275_
timestamp 1644511149
transform 1 0 19504 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1276_
timestamp 1644511149
transform 1 0 33580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1644511149
transform 1 0 2392 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1278_
timestamp 1644511149
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1644511149
transform 1 0 32476 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 1644511149
transform 1 0 25116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1281_
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1644511149
transform 1 0 48116 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1283_
timestamp 1644511149
transform 1 0 30360 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1644511149
transform 1 0 56948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1644511149
transform 1 0 56948 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1644511149
transform 1 0 37996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1287_
timestamp 1644511149
transform 1 0 27968 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1644511149
transform 1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 1644511149
transform 1 0 33120 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 1644511149
transform 1 0 32292 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1292_
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1293_
timestamp 1644511149
transform 1 0 28152 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1295_
timestamp 1644511149
transform 1 0 57132 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1296_
timestamp 1644511149
transform 1 0 57868 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1299_
timestamp 1644511149
transform 1 0 28152 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1644511149
transform 1 0 56948 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 1644511149
transform 1 0 36156 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1644511149
transform 1 0 56488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1305_
timestamp 1644511149
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1306_
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1307_
timestamp 1644511149
transform 1 0 2484 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25944 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31648 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31280 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _1312_
timestamp 1644511149
transform 1 0 28980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1315_
timestamp 1644511149
transform 1 0 30636 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1318_
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1319_
timestamp 1644511149
transform 1 0 28336 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1644511149
transform 1 0 29900 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31464 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31188 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29256 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1324_
timestamp 1644511149
transform 1 0 29716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32476 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1326_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30176 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp 1644511149
transform 1 0 27968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1328_
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1331_
timestamp 1644511149
transform 1 0 31188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1332_
timestamp 1644511149
transform 1 0 29624 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1333_
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1334_
timestamp 1644511149
transform 1 0 33396 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1335_
timestamp 1644511149
transform 1 0 33028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32568 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1337_
timestamp 1644511149
transform 1 0 28612 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _1338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29808 0 1 27200
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_1  _1339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1341_
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30912 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1344_
timestamp 1644511149
transform 1 0 33120 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1345_
timestamp 1644511149
transform 1 0 31556 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1346_
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1347_
timestamp 1644511149
transform 1 0 32384 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1348_
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1349_
timestamp 1644511149
transform 1 0 29624 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30176 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1352_
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1353_
timestamp 1644511149
transform 1 0 31464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1354_
timestamp 1644511149
transform 1 0 29624 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29440 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1356_
timestamp 1644511149
transform 1 0 30728 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1357_
timestamp 1644511149
transform 1 0 29900 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1644511149
transform 1 0 29900 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1359_
timestamp 1644511149
transform 1 0 30268 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1360_
timestamp 1644511149
transform 1 0 29624 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1361_
timestamp 1644511149
transform 1 0 30544 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1362_
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30452 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 1644511149
transform 1 0 33488 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1365_
timestamp 1644511149
transform 1 0 31096 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1366_
timestamp 1644511149
transform 1 0 29900 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1367_
timestamp 1644511149
transform 1 0 28520 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1369_
timestamp 1644511149
transform 1 0 30544 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1370_
timestamp 1644511149
transform 1 0 25484 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1371_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1373_
timestamp 1644511149
transform 1 0 27324 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1374_
timestamp 1644511149
transform 1 0 26128 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1375_
timestamp 1644511149
transform 1 0 29808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1376_
timestamp 1644511149
transform 1 0 26220 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1377_
timestamp 1644511149
transform 1 0 24748 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1379_
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1380_
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1382_
timestamp 1644511149
transform 1 0 25024 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1383_
timestamp 1644511149
transform 1 0 23920 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1384_
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1385_
timestamp 1644511149
transform 1 0 26220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1386_
timestamp 1644511149
transform 1 0 28152 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1387_
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1388_
timestamp 1644511149
transform 1 0 27968 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1389_
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1390_
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1391_
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1392_
timestamp 1644511149
transform 1 0 27508 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1393_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1394_
timestamp 1644511149
transform 1 0 28612 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1396_
timestamp 1644511149
transform 1 0 30820 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1397_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1398_
timestamp 1644511149
transform 1 0 30176 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1399_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1400_
timestamp 1644511149
transform 1 0 30268 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1644511149
transform 1 0 32936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1402_
timestamp 1644511149
transform 1 0 24748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1403_
timestamp 1644511149
transform 1 0 27508 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1404_
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 1644511149
transform 1 0 26036 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1406_
timestamp 1644511149
transform 1 0 24196 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1407_
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1408_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1409_
timestamp 1644511149
transform 1 0 24564 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1410_
timestamp 1644511149
transform 1 0 23552 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1411_
timestamp 1644511149
transform 1 0 24564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1412_
timestamp 1644511149
transform 1 0 23552 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1413_
timestamp 1644511149
transform 1 0 23092 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1644511149
transform 1 0 23736 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1415_
timestamp 1644511149
transform 1 0 24472 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1416_
timestamp 1644511149
transform 1 0 23092 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1418_
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1419_
timestamp 1644511149
transform 1 0 19504 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1420_
timestamp 1644511149
transform 1 0 20976 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1421_
timestamp 1644511149
transform 1 0 27784 0 1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1422_
timestamp 1644511149
transform 1 0 26956 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1423_
timestamp 1644511149
transform 1 0 21252 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1424_
timestamp 1644511149
transform 1 0 22172 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1425_
timestamp 1644511149
transform 1 0 22172 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1426_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1427_
timestamp 1644511149
transform 1 0 20056 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1428_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1429_
timestamp 1644511149
transform 1 0 21712 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1430_
timestamp 1644511149
transform 1 0 20148 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1431_
timestamp 1644511149
transform 1 0 27140 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1433_
timestamp 1644511149
transform 1 0 23920 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1434_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24932 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1435_
timestamp 1644511149
transform 1 0 25944 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1436_
timestamp 1644511149
transform 1 0 25760 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1437_
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1438_
timestamp 1644511149
transform 1 0 22724 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1644511149
transform 1 0 25300 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1440_
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1441_
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1442_
timestamp 1644511149
transform 1 0 23368 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1443_
timestamp 1644511149
transform 1 0 23920 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1444_
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1445_
timestamp 1644511149
transform 1 0 23184 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1446_
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1447_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1448_
timestamp 1644511149
transform 1 0 22724 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1449_
timestamp 1644511149
transform 1 0 22724 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1450_
timestamp 1644511149
transform 1 0 21620 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1451_
timestamp 1644511149
transform 1 0 20976 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1452_
timestamp 1644511149
transform 1 0 19872 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1453_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1454_
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1455_
timestamp 1644511149
transform 1 0 20148 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1456_
timestamp 1644511149
transform 1 0 20884 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1457_
timestamp 1644511149
transform 1 0 20608 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1458_
timestamp 1644511149
transform 1 0 23092 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1459_
timestamp 1644511149
transform 1 0 22816 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1460_
timestamp 1644511149
transform 1 0 24564 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1462_
timestamp 1644511149
transform 1 0 25300 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1644511149
transform 1 0 26128 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1464_
timestamp 1644511149
transform 1 0 25300 0 1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1465_
timestamp 1644511149
transform 1 0 27324 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1466_
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1467_
timestamp 1644511149
transform 1 0 27324 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1468_
timestamp 1644511149
transform 1 0 28428 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1644511149
transform 1 0 27784 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1470_
timestamp 1644511149
transform 1 0 30084 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1471_
timestamp 1644511149
transform 1 0 30912 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1472_
timestamp 1644511149
transform 1 0 29256 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1473_
timestamp 1644511149
transform 1 0 28796 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1474_
timestamp 1644511149
transform 1 0 25392 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1475_
timestamp 1644511149
transform 1 0 29716 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1476_
timestamp 1644511149
transform 1 0 30544 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1477_
timestamp 1644511149
transform 1 0 32108 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1644511149
transform 1 0 32936 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1479_
timestamp 1644511149
transform 1 0 31188 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1644511149
transform 1 0 33856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1481_
timestamp 1644511149
transform 1 0 31188 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 1644511149
transform 1 0 33120 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1483_
timestamp 1644511149
transform 1 0 23644 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1644511149
transform 1 0 22632 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1485_
timestamp 1644511149
transform 1 0 20792 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1644511149
transform 1 0 22540 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1487_
timestamp 1644511149
transform 1 0 23644 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1488_
timestamp 1644511149
transform 1 0 23276 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1644511149
transform 1 0 24748 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1490_
timestamp 1644511149
transform 1 0 22264 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1491_
timestamp 1644511149
transform 1 0 21436 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1492_
timestamp 1644511149
transform 1 0 22540 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1493_
timestamp 1644511149
transform 1 0 21620 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1494_
timestamp 1644511149
transform 1 0 22448 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1495_
timestamp 1644511149
transform 1 0 22172 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1496_
timestamp 1644511149
transform 1 0 23460 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1497_
timestamp 1644511149
transform 1 0 22448 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1498_
timestamp 1644511149
transform 1 0 23276 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1499_
timestamp 1644511149
transform 1 0 23644 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1500_
timestamp 1644511149
transform 1 0 25852 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1501_
timestamp 1644511149
transform 1 0 26220 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1503_
timestamp 1644511149
transform 1 0 27784 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1644511149
transform 1 0 29624 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1505_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1506_
timestamp 1644511149
transform 1 0 27232 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1508_
timestamp 1644511149
transform 1 0 28060 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1509_
timestamp 1644511149
transform 1 0 28336 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1510_
timestamp 1644511149
transform 1 0 28612 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1511_
timestamp 1644511149
transform 1 0 21804 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1644511149
transform 1 0 22356 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1513_
timestamp 1644511149
transform 1 0 26956 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1514_
timestamp 1644511149
transform 1 0 27048 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1515_
timestamp 1644511149
transform 1 0 26036 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1516_
timestamp 1644511149
transform 1 0 29256 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1517_
timestamp 1644511149
transform 1 0 26036 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1518_
timestamp 1644511149
transform 1 0 25392 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1519_
timestamp 1644511149
transform 1 0 25852 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1520_
timestamp 1644511149
transform 1 0 25392 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1521_
timestamp 1644511149
transform 1 0 25392 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1522_
timestamp 1644511149
transform 1 0 26036 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1523_
timestamp 1644511149
transform 1 0 26956 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1524_
timestamp 1644511149
transform 1 0 25576 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1644511149
transform 1 0 27876 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1526_
timestamp 1644511149
transform 1 0 32108 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1527_
timestamp 1644511149
transform 1 0 30360 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1528_
timestamp 1644511149
transform 1 0 33948 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1529_
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1530_
timestamp 1644511149
transform 1 0 29532 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1531_
timestamp 1644511149
transform 1 0 30636 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1532_
timestamp 1644511149
transform 1 0 21712 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1533_
timestamp 1644511149
transform 1 0 21068 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1534_
timestamp 1644511149
transform 1 0 19872 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1535_
timestamp 1644511149
transform 1 0 19228 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1536_
timestamp 1644511149
transform 1 0 19688 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1537_
timestamp 1644511149
transform 1 0 18492 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1538_
timestamp 1644511149
transform 1 0 19412 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1539_
timestamp 1644511149
transform 1 0 18768 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1540_
timestamp 1644511149
transform 1 0 27416 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1541_
timestamp 1644511149
transform 1 0 19596 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1644511149
transform 1 0 20608 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1543_
timestamp 1644511149
transform 1 0 19504 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1544_
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1545_
timestamp 1644511149
transform 1 0 18308 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1546_
timestamp 1644511149
transform 1 0 21068 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1547_
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1548_
timestamp 1644511149
transform 1 0 19504 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1549_
timestamp 1644511149
transform 1 0 26864 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1550_
timestamp 1644511149
transform 1 0 24104 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1551_
timestamp 1644511149
transform 1 0 23736 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1552_
timestamp 1644511149
transform 1 0 23092 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1553_
timestamp 1644511149
transform 1 0 24012 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1556_
timestamp 1644511149
transform 1 0 27784 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1557_
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1558_
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1559_
timestamp 1644511149
transform 1 0 28060 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1560_
timestamp 1644511149
transform 1 0 28152 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1561_
timestamp 1644511149
transform 1 0 27508 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1562_
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1563_
timestamp 1644511149
transform 1 0 20240 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1564_
timestamp 1644511149
transform 1 0 20148 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1565_
timestamp 1644511149
transform 1 0 20056 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1566_
timestamp 1644511149
transform 1 0 21160 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1567_
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1568_
timestamp 1644511149
transform 1 0 32384 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31556 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33672 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1644511149
transform 1 0 29808 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1572_
timestamp 1644511149
transform 1 0 30728 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1573_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1574_
timestamp 1644511149
transform 1 0 31924 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1575_
timestamp 1644511149
transform 1 0 31188 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1576_
timestamp 1644511149
transform 1 0 33948 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1577_
timestamp 1644511149
transform 1 0 33212 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32844 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1579_
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1580_
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1581_
timestamp 1644511149
transform 1 0 25760 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1582_
timestamp 1644511149
transform 1 0 32384 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1583_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1584_
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1585_
timestamp 1644511149
transform 1 0 28244 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1586_
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1587_
timestamp 1644511149
transform 1 0 30636 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1588_
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1589_
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1590_
timestamp 1644511149
transform 1 0 33120 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1591_
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1592_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1593_
timestamp 1644511149
transform 1 0 33028 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1594_
timestamp 1644511149
transform 1 0 31372 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1595_
timestamp 1644511149
transform 1 0 31924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1596_
timestamp 1644511149
transform 1 0 30820 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1597_
timestamp 1644511149
transform 1 0 33028 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1598_
timestamp 1644511149
transform 1 0 36156 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1599_
timestamp 1644511149
transform 1 0 35788 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1600_
timestamp 1644511149
transform 1 0 34132 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1601_
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1602_
timestamp 1644511149
transform 1 0 36708 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1603_
timestamp 1644511149
transform 1 0 40388 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1604_
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1605_
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1606_
timestamp 1644511149
transform 1 0 48668 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1607_
timestamp 1644511149
transform 1 0 47932 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1608_
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1609_
timestamp 1644511149
transform 1 0 33672 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1610_
timestamp 1644511149
transform 1 0 36524 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1611_
timestamp 1644511149
transform 1 0 36432 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1612_
timestamp 1644511149
transform 1 0 39376 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1613_
timestamp 1644511149
transform 1 0 50048 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1614_
timestamp 1644511149
transform 1 0 50508 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1615_
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1616_
timestamp 1644511149
transform 1 0 46736 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1617_
timestamp 1644511149
transform 1 0 37444 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1618_
timestamp 1644511149
transform 1 0 38732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1619_
timestamp 1644511149
transform 1 0 40940 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1620_
timestamp 1644511149
transform 1 0 51428 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1621_
timestamp 1644511149
transform 1 0 53360 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1622_
timestamp 1644511149
transform 1 0 50508 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1623_
timestamp 1644511149
transform 1 0 50508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1624_
timestamp 1644511149
transform 1 0 46736 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1644511149
transform 1 0 36156 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1626_
timestamp 1644511149
transform 1 0 42228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1627_
timestamp 1644511149
transform 1 0 45356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1628_
timestamp 1644511149
transform 1 0 52348 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1629_
timestamp 1644511149
transform 1 0 46736 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1630_
timestamp 1644511149
transform 1 0 38548 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1631_
timestamp 1644511149
transform 1 0 40848 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1632_
timestamp 1644511149
transform 1 0 44068 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1633_
timestamp 1644511149
transform 1 0 50876 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1634_
timestamp 1644511149
transform 1 0 49312 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1636_
timestamp 1644511149
transform 1 0 49220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1637_
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1638_
timestamp 1644511149
transform 1 0 50876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1639_
timestamp 1644511149
transform 1 0 38272 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1640_
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1641_
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1642_
timestamp 1644511149
transform 1 0 42596 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1643_
timestamp 1644511149
transform 1 0 40756 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1644_
timestamp 1644511149
transform 1 0 37812 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1645_
timestamp 1644511149
transform 1 0 49036 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1646_
timestamp 1644511149
transform 1 0 47380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1647_
timestamp 1644511149
transform 1 0 41400 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 1644511149
transform 1 0 36156 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1649_
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1650_
timestamp 1644511149
transform 1 0 31924 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1651_
timestamp 1644511149
transform 1 0 36708 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1652_
timestamp 1644511149
transform 1 0 39376 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1653_
timestamp 1644511149
transform 1 0 37720 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1654_
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1655_
timestamp 1644511149
transform 1 0 40480 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1656_
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1657_
timestamp 1644511149
transform 1 0 34500 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1658_
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1659_
timestamp 1644511149
transform 1 0 49680 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1660_
timestamp 1644511149
transform 1 0 50508 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1661_
timestamp 1644511149
transform 1 0 48392 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1662_
timestamp 1644511149
transform 1 0 34500 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1663_
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1664_
timestamp 1644511149
transform 1 0 50600 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1644511149
transform 1 0 49312 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1666_
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1667_
timestamp 1644511149
transform 1 0 33304 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1668_
timestamp 1644511149
transform 1 0 35696 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1669_
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1670_
timestamp 1644511149
transform 1 0 48116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1671_
timestamp 1644511149
transform 1 0 47932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1672_
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1673_
timestamp 1644511149
transform 1 0 34040 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1674_
timestamp 1644511149
transform 1 0 47840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1675_
timestamp 1644511149
transform 1 0 47932 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1676_
timestamp 1644511149
transform 1 0 33396 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1677_
timestamp 1644511149
transform 1 0 32200 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1678_
timestamp 1644511149
transform 1 0 49680 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1679_
timestamp 1644511149
transform 1 0 51888 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1680_
timestamp 1644511149
transform 1 0 42780 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1681_
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1682_
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1683_
timestamp 1644511149
transform 1 0 35696 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1684_
timestamp 1644511149
transform 1 0 36616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1685_
timestamp 1644511149
transform 1 0 35696 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1686_
timestamp 1644511149
transform 1 0 35052 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1687_
timestamp 1644511149
transform 1 0 37536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1688_
timestamp 1644511149
transform 1 0 41216 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1689_
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1690_
timestamp 1644511149
transform 1 0 35144 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1691_
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1692_
timestamp 1644511149
transform 1 0 35696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1693_
timestamp 1644511149
transform 1 0 35328 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1694_
timestamp 1644511149
transform 1 0 34132 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1695_
timestamp 1644511149
transform 1 0 27140 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1696_
timestamp 1644511149
transform 1 0 35512 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1697_
timestamp 1644511149
transform 1 0 40664 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1698_
timestamp 1644511149
transform 1 0 39376 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1699_
timestamp 1644511149
transform 1 0 38916 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1700_
timestamp 1644511149
transform 1 0 40756 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1701_
timestamp 1644511149
transform 1 0 40388 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1702_
timestamp 1644511149
transform 1 0 39928 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1703_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38272 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1704_
timestamp 1644511149
transform 1 0 39284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1705_
timestamp 1644511149
transform 1 0 37444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1706_
timestamp 1644511149
transform 1 0 36064 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1707_
timestamp 1644511149
transform 1 0 36616 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1708_
timestamp 1644511149
transform 1 0 36432 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1709_
timestamp 1644511149
transform 1 0 39928 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1710_
timestamp 1644511149
transform 1 0 38824 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1711_
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1712_
timestamp 1644511149
transform 1 0 36156 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36800 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1714_
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1715_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36340 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1716_
timestamp 1644511149
transform 1 0 38548 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1717_
timestamp 1644511149
transform 1 0 39192 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1718_
timestamp 1644511149
transform 1 0 37720 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38548 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1720_
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_4  _1721_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _1722_
timestamp 1644511149
transform 1 0 37352 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1723_
timestamp 1644511149
transform 1 0 36248 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1724_
timestamp 1644511149
transform 1 0 37260 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1725_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1726_
timestamp 1644511149
transform 1 0 40848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1727_
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _1728_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1729_
timestamp 1644511149
transform 1 0 37352 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1730_
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1731_
timestamp 1644511149
transform 1 0 40204 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1732_
timestamp 1644511149
transform 1 0 40112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1733_
timestamp 1644511149
transform 1 0 38548 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1734_
timestamp 1644511149
transform 1 0 38456 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1735_
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _1736_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40848 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1737_
timestamp 1644511149
transform 1 0 41676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1738_
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1739_
timestamp 1644511149
transform 1 0 37536 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1740_
timestamp 1644511149
transform 1 0 39560 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1741_
timestamp 1644511149
transform 1 0 41400 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1742_
timestamp 1644511149
transform 1 0 43332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1743_
timestamp 1644511149
transform 1 0 42596 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1744_
timestamp 1644511149
transform 1 0 38272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1745_
timestamp 1644511149
transform 1 0 39192 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1746_
timestamp 1644511149
transform 1 0 39928 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1747_
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1748_
timestamp 1644511149
transform 1 0 41032 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1749_
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1750_
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1751_
timestamp 1644511149
transform 1 0 38916 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1752_
timestamp 1644511149
transform 1 0 41860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1753_
timestamp 1644511149
transform 1 0 40664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1754_
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1755_
timestamp 1644511149
transform 1 0 40848 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1756_
timestamp 1644511149
transform 1 0 42780 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1757_
timestamp 1644511149
transform 1 0 43332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1758_
timestamp 1644511149
transform 1 0 48852 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1759_
timestamp 1644511149
transform 1 0 47748 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1761_
timestamp 1644511149
transform 1 0 41400 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1762_
timestamp 1644511149
transform 1 0 46276 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1644511149
transform 1 0 47104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1764_
timestamp 1644511149
transform 1 0 46368 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1765_
timestamp 1644511149
transform 1 0 44160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1766_
timestamp 1644511149
transform 1 0 45172 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1767_
timestamp 1644511149
transform 1 0 42412 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1768_
timestamp 1644511149
transform 1 0 43056 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1769_
timestamp 1644511149
transform 1 0 43424 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1770_
timestamp 1644511149
transform 1 0 45264 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1771_
timestamp 1644511149
transform 1 0 43884 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1772_
timestamp 1644511149
transform 1 0 44068 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1773_
timestamp 1644511149
transform 1 0 41400 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1774_
timestamp 1644511149
transform 1 0 43700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1775_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44252 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1776_
timestamp 1644511149
transform 1 0 41308 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1777_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46276 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1644511149
transform 1 0 44068 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1779_
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1780_
timestamp 1644511149
transform 1 0 43424 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _1781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43240 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1782_
timestamp 1644511149
transform 1 0 43332 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1783_
timestamp 1644511149
transform 1 0 44068 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1784_
timestamp 1644511149
transform 1 0 43332 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1785_
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1786_
timestamp 1644511149
transform 1 0 44160 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1788_
timestamp 1644511149
transform 1 0 43148 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1789_
timestamp 1644511149
transform 1 0 44804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1790_
timestamp 1644511149
transform 1 0 45816 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1791_
timestamp 1644511149
transform 1 0 48852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1792_
timestamp 1644511149
transform 1 0 46920 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1793_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1794_
timestamp 1644511149
transform 1 0 47840 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 1644511149
transform 1 0 46644 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1796_
timestamp 1644511149
transform 1 0 46460 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1797_
timestamp 1644511149
transform 1 0 48024 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1798_
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1799_
timestamp 1644511149
transform 1 0 49404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1800_
timestamp 1644511149
transform 1 0 48852 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1801_
timestamp 1644511149
transform 1 0 47932 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1802_
timestamp 1644511149
transform 1 0 47104 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1803_
timestamp 1644511149
transform 1 0 47380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1804_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1805_
timestamp 1644511149
transform 1 0 46460 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1806_
timestamp 1644511149
transform 1 0 45908 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1807_
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1808_
timestamp 1644511149
transform 1 0 44068 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1809_
timestamp 1644511149
transform 1 0 43792 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1810_
timestamp 1644511149
transform 1 0 44160 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_1  _1811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43148 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1812_
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1813_
timestamp 1644511149
transform 1 0 45448 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1814_
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1815_
timestamp 1644511149
transform 1 0 44988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1816_
timestamp 1644511149
transform 1 0 44804 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1817_
timestamp 1644511149
transform 1 0 43424 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1818_
timestamp 1644511149
transform 1 0 42504 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1819_
timestamp 1644511149
transform 1 0 41860 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1820_
timestamp 1644511149
transform 1 0 43240 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1821_
timestamp 1644511149
transform 1 0 41768 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1823_
timestamp 1644511149
transform 1 0 41676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1824_
timestamp 1644511149
transform 1 0 43424 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1825_
timestamp 1644511149
transform 1 0 45264 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1826_
timestamp 1644511149
transform 1 0 44804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1827_
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1828_
timestamp 1644511149
transform 1 0 43608 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1829_
timestamp 1644511149
transform 1 0 43700 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1830_
timestamp 1644511149
transform 1 0 43792 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1831_
timestamp 1644511149
transform 1 0 44068 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1832_
timestamp 1644511149
transform 1 0 43884 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1833_
timestamp 1644511149
transform 1 0 46276 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1834_
timestamp 1644511149
transform 1 0 45908 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1835_
timestamp 1644511149
transform 1 0 45448 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1836_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46092 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1837_
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1838_
timestamp 1644511149
transform 1 0 45816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1839_
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1840_
timestamp 1644511149
transform 1 0 47380 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1841_
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1842_
timestamp 1644511149
transform 1 0 46368 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1843_
timestamp 1644511149
transform 1 0 41124 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1844_
timestamp 1644511149
transform 1 0 47104 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1845_
timestamp 1644511149
transform 1 0 50600 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1846_
timestamp 1644511149
transform 1 0 50784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1847_
timestamp 1644511149
transform 1 0 47012 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1848_
timestamp 1644511149
transform 1 0 49956 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1849_
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1850_
timestamp 1644511149
transform 1 0 47656 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1851_
timestamp 1644511149
transform 1 0 46276 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1852_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1853_
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1854_
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1855_
timestamp 1644511149
transform 1 0 48024 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1856_
timestamp 1644511149
transform 1 0 46460 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1857_
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1858_
timestamp 1644511149
transform 1 0 44068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1859_
timestamp 1644511149
transform 1 0 42780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1860_
timestamp 1644511149
transform 1 0 44712 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1861_
timestamp 1644511149
transform 1 0 42964 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1862_
timestamp 1644511149
transform 1 0 40204 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1863_
timestamp 1644511149
transform 1 0 42688 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1864_
timestamp 1644511149
transform 1 0 42320 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _1865_
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 1644511149
transform 1 0 41492 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1867_
timestamp 1644511149
transform 1 0 41308 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1868_
timestamp 1644511149
transform 1 0 40940 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1869_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43884 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1870_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1871_
timestamp 1644511149
transform 1 0 44896 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1872_
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1873_
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _1874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43608 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1875_
timestamp 1644511149
transform 1 0 45908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1876_
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1877_
timestamp 1644511149
transform 1 0 44068 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1878_
timestamp 1644511149
transform 1 0 40480 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1879_
timestamp 1644511149
transform 1 0 41032 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1880_
timestamp 1644511149
transform 1 0 41492 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1881_
timestamp 1644511149
transform 1 0 41492 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1882_
timestamp 1644511149
transform 1 0 40296 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1883_
timestamp 1644511149
transform 1 0 39928 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1884_
timestamp 1644511149
transform 1 0 45448 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1885_
timestamp 1644511149
transform 1 0 43424 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1886_
timestamp 1644511149
transform 1 0 43976 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1887_
timestamp 1644511149
transform 1 0 42964 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1888_
timestamp 1644511149
transform 1 0 42964 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1889_
timestamp 1644511149
transform 1 0 44252 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1890_
timestamp 1644511149
transform 1 0 45080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _1891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43516 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1892_
timestamp 1644511149
transform 1 0 41216 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1893_
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1894_
timestamp 1644511149
transform 1 0 46460 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1895_
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46736 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2oi_1  _1897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48024 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1898_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45540 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1899_
timestamp 1644511149
transform 1 0 45632 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1900_
timestamp 1644511149
transform 1 0 47104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1901_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1902_
timestamp 1644511149
transform 1 0 47840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1903_
timestamp 1644511149
transform 1 0 47012 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1904_
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1905_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1906_
timestamp 1644511149
transform 1 0 44068 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1907_
timestamp 1644511149
transform 1 0 50692 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1908_
timestamp 1644511149
transform 1 0 49128 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1909_
timestamp 1644511149
transform 1 0 44896 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1910_
timestamp 1644511149
transform 1 0 43424 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1911_
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1912_
timestamp 1644511149
transform 1 0 44436 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1913_
timestamp 1644511149
transform 1 0 44436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1914_
timestamp 1644511149
transform 1 0 43608 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1915_
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1916_
timestamp 1644511149
transform 1 0 44436 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1917_
timestamp 1644511149
transform 1 0 43240 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1918_
timestamp 1644511149
transform 1 0 40572 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1919_
timestamp 1644511149
transform 1 0 41308 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1920_
timestamp 1644511149
transform 1 0 40388 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1921_
timestamp 1644511149
transform 1 0 41676 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1922_
timestamp 1644511149
transform 1 0 42044 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_2  _1923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1924_
timestamp 1644511149
transform 1 0 47656 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1925_
timestamp 1644511149
transform 1 0 43608 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _1926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42044 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1927_
timestamp 1644511149
transform 1 0 45356 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1928_
timestamp 1644511149
transform 1 0 40112 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1930_
timestamp 1644511149
transform 1 0 41124 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1931_
timestamp 1644511149
transform 1 0 43976 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _1932_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39192 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1933_
timestamp 1644511149
transform 1 0 53084 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1934_
timestamp 1644511149
transform 1 0 48484 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1935_
timestamp 1644511149
transform 1 0 44344 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1936_
timestamp 1644511149
transform 1 0 39560 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1937_
timestamp 1644511149
transform 1 0 41308 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _1938_
timestamp 1644511149
transform 1 0 40572 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1939_
timestamp 1644511149
transform 1 0 44068 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1940_
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _1941_
timestamp 1644511149
transform 1 0 43608 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1942_
timestamp 1644511149
transform 1 0 29992 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1943_
timestamp 1644511149
transform 1 0 34776 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1944_
timestamp 1644511149
transform 1 0 42872 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1945_
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1946_
timestamp 1644511149
transform 1 0 49036 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1947_
timestamp 1644511149
transform 1 0 48852 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1948_
timestamp 1644511149
transform 1 0 47104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1949_
timestamp 1644511149
transform 1 0 46460 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1950_
timestamp 1644511149
transform 1 0 46736 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _1951_
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1952_
timestamp 1644511149
transform 1 0 45448 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1953_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _1954_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46276 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1955_
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1956_
timestamp 1644511149
transform 1 0 45264 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1957_
timestamp 1644511149
transform 1 0 47196 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1958_
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1959_
timestamp 1644511149
transform 1 0 46460 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1960_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1961_
timestamp 1644511149
transform 1 0 42136 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1962_
timestamp 1644511149
transform 1 0 42964 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1963_
timestamp 1644511149
transform 1 0 45724 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1964_
timestamp 1644511149
transform 1 0 46092 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1965_
timestamp 1644511149
transform 1 0 43884 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1966_
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1967_
timestamp 1644511149
transform 1 0 49956 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1968_
timestamp 1644511149
transform 1 0 51244 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50324 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1970_
timestamp 1644511149
transform 1 0 51428 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50140 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1972_
timestamp 1644511149
transform 1 0 50048 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1973_
timestamp 1644511149
transform 1 0 49128 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1974_
timestamp 1644511149
transform 1 0 49220 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1975_
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1976_
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1977_
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1978_
timestamp 1644511149
transform 1 0 47748 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1979_
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1980_
timestamp 1644511149
transform 1 0 44804 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1981_
timestamp 1644511149
transform 1 0 46828 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1982_
timestamp 1644511149
transform 1 0 41308 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1983_
timestamp 1644511149
transform 1 0 46000 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1984_
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1985_
timestamp 1644511149
transform 1 0 44988 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1986_
timestamp 1644511149
transform 1 0 48300 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1987_
timestamp 1644511149
transform 1 0 47564 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1988_
timestamp 1644511149
transform 1 0 46736 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1989_
timestamp 1644511149
transform 1 0 47656 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1990_
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_2  _1991_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48576 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1992_
timestamp 1644511149
transform 1 0 41952 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1993_
timestamp 1644511149
transform 1 0 32568 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1994_
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1995_
timestamp 1644511149
transform 1 0 50140 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1996_
timestamp 1644511149
transform 1 0 50784 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1997_
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1998_
timestamp 1644511149
transform 1 0 45632 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1999_
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2000_
timestamp 1644511149
transform 1 0 42688 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2001_
timestamp 1644511149
transform 1 0 43332 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2002_
timestamp 1644511149
transform 1 0 50784 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2003_
timestamp 1644511149
transform 1 0 50140 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2004_
timestamp 1644511149
transform 1 0 50784 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2005_
timestamp 1644511149
transform 1 0 51796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2006_
timestamp 1644511149
transform 1 0 51796 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2007_
timestamp 1644511149
transform 1 0 49956 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2008_
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2009_
timestamp 1644511149
transform 1 0 51244 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2010_
timestamp 1644511149
transform 1 0 50508 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2011_
timestamp 1644511149
transform 1 0 48116 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2012_
timestamp 1644511149
transform 1 0 49864 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2013_
timestamp 1644511149
transform 1 0 50140 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2014_
timestamp 1644511149
transform 1 0 45540 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2015_
timestamp 1644511149
transform 1 0 46828 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2016_
timestamp 1644511149
transform 1 0 49864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2017_
timestamp 1644511149
transform 1 0 47932 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2018_
timestamp 1644511149
transform 1 0 48668 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2019_
timestamp 1644511149
transform 1 0 48668 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2020_
timestamp 1644511149
transform 1 0 44712 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2021_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46092 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2022_
timestamp 1644511149
transform 1 0 44160 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2023_
timestamp 1644511149
transform 1 0 46000 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2024_
timestamp 1644511149
transform 1 0 44712 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2025_
timestamp 1644511149
transform 1 0 35052 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2026_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2027_
timestamp 1644511149
transform 1 0 50784 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _2028_
timestamp 1644511149
transform 1 0 49864 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2029_
timestamp 1644511149
transform 1 0 50968 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2030_
timestamp 1644511149
transform 1 0 51704 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2031_
timestamp 1644511149
transform 1 0 52716 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2032_
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2033_
timestamp 1644511149
transform 1 0 52072 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2034_
timestamp 1644511149
transform 1 0 52256 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2035_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2036_
timestamp 1644511149
transform 1 0 53452 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2037_
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2038_
timestamp 1644511149
transform 1 0 52624 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2039_
timestamp 1644511149
transform 1 0 53084 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2040_
timestamp 1644511149
transform 1 0 52532 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2041_
timestamp 1644511149
transform 1 0 52072 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2042_
timestamp 1644511149
transform 1 0 51980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2043_
timestamp 1644511149
transform 1 0 51428 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2044_
timestamp 1644511149
transform 1 0 42780 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2045_
timestamp 1644511149
transform 1 0 42412 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2046_
timestamp 1644511149
transform 1 0 42872 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2047_
timestamp 1644511149
transform 1 0 44068 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2048_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _2049_
timestamp 1644511149
transform 1 0 42136 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2050_
timestamp 1644511149
transform 1 0 43240 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2051_
timestamp 1644511149
transform 1 0 47472 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2052_
timestamp 1644511149
transform 1 0 47748 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2053_
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _2054_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2055_
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2056_
timestamp 1644511149
transform 1 0 41584 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2057_
timestamp 1644511149
transform 1 0 42412 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2058_
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2059_
timestamp 1644511149
transform 1 0 51152 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2060_
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _2061_
timestamp 1644511149
transform 1 0 42504 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2062_
timestamp 1644511149
transform 1 0 43424 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2063_
timestamp 1644511149
transform 1 0 50508 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2064_
timestamp 1644511149
transform 1 0 35328 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_2  _2065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52716 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _2066_
timestamp 1644511149
transform 1 0 48392 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2067_
timestamp 1644511149
transform 1 0 51244 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2068_
timestamp 1644511149
transform 1 0 53912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2069_
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_1  _2070_
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2071_
timestamp 1644511149
transform 1 0 51060 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _2072_
timestamp 1644511149
transform 1 0 50968 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _2073_
timestamp 1644511149
transform 1 0 51336 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2074_
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2075_
timestamp 1644511149
transform 1 0 53176 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2076_
timestamp 1644511149
transform 1 0 53452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2077_
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2078_
timestamp 1644511149
transform 1 0 53912 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2079_
timestamp 1644511149
transform 1 0 53820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2080_
timestamp 1644511149
transform 1 0 54464 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2081_
timestamp 1644511149
transform 1 0 54188 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2082_
timestamp 1644511149
transform 1 0 54556 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2083_
timestamp 1644511149
transform 1 0 53912 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2084_
timestamp 1644511149
transform 1 0 54188 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2085_
timestamp 1644511149
transform 1 0 54004 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2086_
timestamp 1644511149
transform 1 0 53728 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2087_
timestamp 1644511149
transform 1 0 53544 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2088_
timestamp 1644511149
transform 1 0 52532 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2089_
timestamp 1644511149
transform 1 0 53452 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2090_
timestamp 1644511149
transform 1 0 39192 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2091_
timestamp 1644511149
transform 1 0 37536 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2092_
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2093_
timestamp 1644511149
transform 1 0 37996 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _2094_
timestamp 1644511149
transform 1 0 37628 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2095_
timestamp 1644511149
transform 1 0 38088 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2096_
timestamp 1644511149
transform 1 0 38824 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2097_
timestamp 1644511149
transform 1 0 39100 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2098_
timestamp 1644511149
transform 1 0 38088 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2099_
timestamp 1644511149
transform 1 0 51612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _2100_
timestamp 1644511149
transform 1 0 39928 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2101_
timestamp 1644511149
transform 1 0 39836 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _2102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38732 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2103_
timestamp 1644511149
transform 1 0 37720 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2104_
timestamp 1644511149
transform 1 0 37076 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2105_
timestamp 1644511149
transform 1 0 34960 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2106_
timestamp 1644511149
transform 1 0 48024 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2107_
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2108_
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2109_
timestamp 1644511149
transform 1 0 41492 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2110_
timestamp 1644511149
transform 1 0 40480 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2111_
timestamp 1644511149
transform 1 0 39652 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2112_
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2113_
timestamp 1644511149
transform 1 0 37260 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _2114_
timestamp 1644511149
transform 1 0 54924 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2115_
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2116_
timestamp 1644511149
transform 1 0 55292 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2117_
timestamp 1644511149
transform 1 0 41216 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2118_
timestamp 1644511149
transform 1 0 51428 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2119_
timestamp 1644511149
transform 1 0 55200 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2120_
timestamp 1644511149
transform 1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2121_
timestamp 1644511149
transform 1 0 51336 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2122_
timestamp 1644511149
transform 1 0 49496 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2123_
timestamp 1644511149
transform 1 0 51520 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2124_
timestamp 1644511149
transform 1 0 51428 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2125_
timestamp 1644511149
transform 1 0 50600 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2126_
timestamp 1644511149
transform 1 0 49036 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _2127_
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _2128_
timestamp 1644511149
transform 1 0 52716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _2129_
timestamp 1644511149
transform 1 0 52256 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2130_
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2131_
timestamp 1644511149
transform 1 0 54464 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2132_
timestamp 1644511149
transform 1 0 54280 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2133_
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2134_
timestamp 1644511149
transform 1 0 55384 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2135_
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2136_
timestamp 1644511149
transform 1 0 55660 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2137_
timestamp 1644511149
transform 1 0 54740 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2138_
timestamp 1644511149
transform 1 0 55476 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2139_
timestamp 1644511149
transform 1 0 55476 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2140_
timestamp 1644511149
transform 1 0 55844 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2141_
timestamp 1644511149
transform 1 0 55936 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2142_
timestamp 1644511149
transform 1 0 57132 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2143_
timestamp 1644511149
transform 1 0 56304 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2144_
timestamp 1644511149
transform 1 0 56212 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2145_
timestamp 1644511149
transform 1 0 55108 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2146_
timestamp 1644511149
transform 1 0 55292 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2147_
timestamp 1644511149
transform 1 0 54464 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2148_
timestamp 1644511149
transform 1 0 55292 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2149_
timestamp 1644511149
transform 1 0 54372 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2150_
timestamp 1644511149
transform 1 0 38456 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2151_
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2152_
timestamp 1644511149
transform 1 0 41124 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2153_
timestamp 1644511149
transform 1 0 41308 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _2154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40940 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _2155_
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2156_
timestamp 1644511149
transform 1 0 37904 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2157_
timestamp 1644511149
transform 1 0 36432 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2158_
timestamp 1644511149
transform 1 0 37352 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2159_
timestamp 1644511149
transform 1 0 35972 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2160_
timestamp 1644511149
transform 1 0 35972 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2161_
timestamp 1644511149
transform 1 0 40940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _2162_
timestamp 1644511149
transform 1 0 41400 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2163_
timestamp 1644511149
transform 1 0 41032 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2164_
timestamp 1644511149
transform 1 0 42136 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2165_
timestamp 1644511149
transform 1 0 39560 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2166_
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2167_
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _2168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40204 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2169_
timestamp 1644511149
transform 1 0 55200 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _2170_
timestamp 1644511149
transform 1 0 56304 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2171_
timestamp 1644511149
transform 1 0 56120 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2172_
timestamp 1644511149
transform 1 0 56212 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2173_
timestamp 1644511149
transform 1 0 52624 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2174_
timestamp 1644511149
transform 1 0 51428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2175_
timestamp 1644511149
transform 1 0 51796 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2176_
timestamp 1644511149
transform 1 0 53176 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2177_
timestamp 1644511149
transform 1 0 53360 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2178_
timestamp 1644511149
transform 1 0 49036 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2179_
timestamp 1644511149
transform 1 0 50508 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2180_
timestamp 1644511149
transform 1 0 50416 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2181_
timestamp 1644511149
transform 1 0 50876 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2182_
timestamp 1644511149
transform 1 0 51704 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2183_
timestamp 1644511149
transform 1 0 51796 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2184_
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2185_
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2186_
timestamp 1644511149
transform 1 0 49404 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2187_
timestamp 1644511149
transform 1 0 49128 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _2188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48852 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2189_
timestamp 1644511149
transform 1 0 52624 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2190_
timestamp 1644511149
transform 1 0 53912 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2191_
timestamp 1644511149
transform 1 0 54464 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2192_
timestamp 1644511149
transform 1 0 54556 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2193_
timestamp 1644511149
transform 1 0 55384 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2194_
timestamp 1644511149
transform 1 0 55568 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2195_
timestamp 1644511149
transform 1 0 56488 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2196_
timestamp 1644511149
transform 1 0 55476 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2197_
timestamp 1644511149
transform 1 0 56304 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2198_
timestamp 1644511149
transform 1 0 56948 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2199_
timestamp 1644511149
transform 1 0 56856 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2200_
timestamp 1644511149
transform 1 0 56856 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2201_
timestamp 1644511149
transform 1 0 56856 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2202_
timestamp 1644511149
transform 1 0 56580 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2203_
timestamp 1644511149
transform 1 0 56672 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2204_
timestamp 1644511149
transform 1 0 56856 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2205_
timestamp 1644511149
transform 1 0 56856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _2206_
timestamp 1644511149
transform 1 0 56028 0 -1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _2207_
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2208_
timestamp 1644511149
transform 1 0 40480 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2209_
timestamp 1644511149
transform 1 0 36984 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2210_
timestamp 1644511149
transform 1 0 37076 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2211_
timestamp 1644511149
transform 1 0 38272 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2212_
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2213_
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2214_
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2215_
timestamp 1644511149
transform 1 0 38548 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2216_
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2217_
timestamp 1644511149
transform 1 0 33120 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2218_
timestamp 1644511149
transform 1 0 56304 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2219_
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2220_
timestamp 1644511149
transform 1 0 57776 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _2221_
timestamp 1644511149
transform 1 0 55844 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2222_
timestamp 1644511149
transform 1 0 54004 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2223_
timestamp 1644511149
transform 1 0 48576 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2224_
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2225_
timestamp 1644511149
transform 1 0 51980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2226_
timestamp 1644511149
transform 1 0 51336 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2227_
timestamp 1644511149
transform 1 0 50600 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2228_
timestamp 1644511149
transform 1 0 52716 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2229_
timestamp 1644511149
transform 1 0 52900 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2230_
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2231_
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2232_
timestamp 1644511149
transform 1 0 50692 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2233_
timestamp 1644511149
transform 1 0 52164 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2234_
timestamp 1644511149
transform 1 0 48852 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2235_
timestamp 1644511149
transform 1 0 48576 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2236_
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2237_
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2238_
timestamp 1644511149
transform 1 0 50600 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2239_
timestamp 1644511149
transform 1 0 52164 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2240_
timestamp 1644511149
transform 1 0 53176 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2241_
timestamp 1644511149
transform 1 0 54832 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2242_
timestamp 1644511149
transform 1 0 55844 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2243_
timestamp 1644511149
transform 1 0 56212 0 1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _2244_
timestamp 1644511149
transform 1 0 55752 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _2245_
timestamp 1644511149
transform 1 0 55292 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2246_
timestamp 1644511149
transform 1 0 41308 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2247_
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2248_
timestamp 1644511149
transform 1 0 41032 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2249_
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2250_
timestamp 1644511149
transform 1 0 38548 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2251_
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _2252_
timestamp 1644511149
transform 1 0 40296 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2253_
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2254_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2255_
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2256_
timestamp 1644511149
transform 1 0 33028 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2258_
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2259_
timestamp 1644511149
transform 1 0 24840 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2260_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2261_
timestamp 1644511149
transform 1 0 27508 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2262_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2263_
timestamp 1644511149
transform 1 0 27600 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2264_
timestamp 1644511149
transform 1 0 31004 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2265_
timestamp 1644511149
transform 1 0 31096 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2266_
timestamp 1644511149
transform 1 0 23828 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2267_
timestamp 1644511149
transform 1 0 21160 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2268_
timestamp 1644511149
transform 1 0 19504 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2269_
timestamp 1644511149
transform 1 0 25300 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2270_
timestamp 1644511149
transform 1 0 24380 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2271_
timestamp 1644511149
transform 1 0 21344 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2272_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2274_
timestamp 1644511149
transform 1 0 27600 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2275_
timestamp 1644511149
transform 1 0 27600 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2276_
timestamp 1644511149
transform 1 0 28244 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2277_
timestamp 1644511149
transform 1 0 28520 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2278_
timestamp 1644511149
transform 1 0 30176 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2279_
timestamp 1644511149
transform 1 0 32016 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2280_
timestamp 1644511149
transform 1 0 32108 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2281_
timestamp 1644511149
transform 1 0 32108 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2282_
timestamp 1644511149
transform 1 0 22356 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2283_
timestamp 1644511149
transform 1 0 21804 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2284_
timestamp 1644511149
transform 1 0 22080 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2285_
timestamp 1644511149
transform 1 0 21896 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2286_
timestamp 1644511149
transform 1 0 21804 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2287_
timestamp 1644511149
transform 1 0 21620 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2288_
timestamp 1644511149
transform 1 0 22080 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2289_
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2290_
timestamp 1644511149
transform 1 0 25024 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2291_
timestamp 1644511149
transform 1 0 29532 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2292_
timestamp 1644511149
transform 1 0 23000 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2293_
timestamp 1644511149
transform 1 0 27048 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2294_
timestamp 1644511149
transform 1 0 29532 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2295_
timestamp 1644511149
transform 1 0 27416 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2296_
timestamp 1644511149
transform 1 0 24932 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2297_
timestamp 1644511149
transform 1 0 25116 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2298_
timestamp 1644511149
transform 1 0 25484 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2299_
timestamp 1644511149
transform 1 0 25024 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2300_
timestamp 1644511149
transform 1 0 27600 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2301_
timestamp 1644511149
transform 1 0 20056 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2302_
timestamp 1644511149
transform 1 0 19228 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2303_
timestamp 1644511149
transform 1 0 19228 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2304_
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2305_
timestamp 1644511149
transform 1 0 18768 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2306_
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2307_
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2308_
timestamp 1644511149
transform 1 0 19044 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2309_
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2310_
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2311_
timestamp 1644511149
transform 1 0 30084 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2312_
timestamp 1644511149
transform 1 0 27600 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2313_
timestamp 1644511149
transform 1 0 21712 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _2314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2315_
timestamp 1644511149
transform 1 0 27876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2316_
timestamp 1644511149
transform 1 0 27600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2317_
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2318_
timestamp 1644511149
transform 1 0 30728 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2319_
timestamp 1644511149
transform 1 0 25024 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2320_
timestamp 1644511149
transform 1 0 24840 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2321_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2322_
timestamp 1644511149
transform 1 0 27508 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2323_
timestamp 1644511149
transform 1 0 27876 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2324_
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2325_
timestamp 1644511149
transform 1 0 30912 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2326_
timestamp 1644511149
transform 1 0 30176 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2327_
timestamp 1644511149
transform 1 0 34132 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2328_
timestamp 1644511149
transform 1 0 34960 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2329_
timestamp 1644511149
transform 1 0 36800 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2330_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2331_
timestamp 1644511149
transform 1 0 37168 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2332_
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2333_
timestamp 1644511149
transform 1 0 37168 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2334_
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2335_
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2336_
timestamp 1644511149
transform 1 0 37352 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2337_
timestamp 1644511149
transform 1 0 37352 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2338_
timestamp 1644511149
transform 1 0 37536 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2339_
timestamp 1644511149
transform 1 0 29992 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2340_
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2341_
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2342_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2343_
timestamp 1644511149
transform 1 0 33856 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2344_
timestamp 1644511149
transform 1 0 33764 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2345_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2346_
timestamp 1644511149
transform 1 0 34132 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2347_
timestamp 1644511149
transform 1 0 34040 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2348_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2349_
timestamp 1644511149
transform 1 0 34224 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2350_
timestamp 1644511149
transform 1 0 31096 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2351_
timestamp 1644511149
transform 1 0 30728 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2352_
timestamp 1644511149
transform 1 0 31004 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2353_
timestamp 1644511149
transform 1 0 33488 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2354_
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2355_
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2356_
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2357_
timestamp 1644511149
transform 1 0 32752 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _2358__7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2359__8
timestamp 1644511149
transform 1 0 2024 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2360__9
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2361__10
timestamp 1644511149
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2362__11
timestamp 1644511149
transform 1 0 54004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2363__12
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2364__13
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2365__14
timestamp 1644511149
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2366__15
timestamp 1644511149
transform 1 0 57868 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2367__16
timestamp 1644511149
transform 1 0 55660 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2368__17
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2369__18
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2370__19
timestamp 1644511149
transform 1 0 57868 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2371__20
timestamp 1644511149
transform 1 0 6256 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2372__21
timestamp 1644511149
transform 1 0 32108 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2373__22
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2374__23
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2375__24
timestamp 1644511149
transform 1 0 57868 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2376__25
timestamp 1644511149
transform 1 0 7452 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2377__26
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2378__27
timestamp 1644511149
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2379__28
timestamp 1644511149
transform 1 0 57592 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2380__29
timestamp 1644511149
transform 1 0 35788 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2381__30
timestamp 1644511149
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2382__31
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2383__32
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2384__33
timestamp 1644511149
transform 1 0 57592 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2385__34
timestamp 1644511149
transform 1 0 2024 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2386__35
timestamp 1644511149
transform 1 0 53360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2387__36
timestamp 1644511149
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2388__37
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2389__38
timestamp 1644511149
transform 1 0 57868 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2390__39
timestamp 1644511149
transform 1 0 56488 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2391__40
timestamp 1644511149
transform 1 0 39836 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2392__41
timestamp 1644511149
transform 1 0 8096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2393__42
timestamp 1644511149
transform 1 0 2944 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2394__43
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2395__44
timestamp 1644511149
transform 1 0 27692 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2396__45
timestamp 1644511149
transform 1 0 55844 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2397__46
timestamp 1644511149
transform 1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2398__47
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2399__48
timestamp 1644511149
transform 1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2400__49
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2401__50
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2402__51
timestamp 1644511149
transform 1 0 38364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2403__52
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2404__53
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2405__54
timestamp 1644511149
transform 1 0 42688 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2406__55
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2407__56
timestamp 1644511149
transform 1 0 46276 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2408__57
timestamp 1644511149
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2409__58
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2410__59
timestamp 1644511149
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2411__60
timestamp 1644511149
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2412__61
timestamp 1644511149
transform 1 0 2668 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2413__62
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2414__63
timestamp 1644511149
transform 1 0 57684 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2415__64
timestamp 1644511149
transform 1 0 57592 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2416__65
timestamp 1644511149
transform 1 0 19228 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2417__66
timestamp 1644511149
transform 1 0 57868 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2418__67
timestamp 1644511149
transform 1 0 30452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2419__68
timestamp 1644511149
transform 1 0 46276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2420__69
timestamp 1644511149
transform 1 0 50140 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2421__70
timestamp 1644511149
transform 1 0 29808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2422__71
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2423__72
timestamp 1644511149
transform 1 0 2208 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2424__73
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2425__74
timestamp 1644511149
transform 1 0 15824 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2426__75
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2427__76
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2428__77
timestamp 1644511149
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2429__78
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2430__79
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2431__80
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2432__81
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2433__82
timestamp 1644511149
transform 1 0 18032 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2434__83
timestamp 1644511149
transform 1 0 55660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2435__84
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2436__85
timestamp 1644511149
transform 1 0 42044 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2437__86
timestamp 1644511149
transform 1 0 17756 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2438__87
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2439__88
timestamp 1644511149
transform 1 0 2668 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2440__89
timestamp 1644511149
transform 1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2441__90
timestamp 1644511149
transform 1 0 29992 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2442__91
timestamp 1644511149
transform 1 0 31280 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2443__92
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2444__93
timestamp 1644511149
transform 1 0 57868 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2445__94
timestamp 1644511149
transform 1 0 35696 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2446__95
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2447__96
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2448__97
timestamp 1644511149
transform 1 0 3864 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2449__98
timestamp 1644511149
transform 1 0 48576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2450__99
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2451__100
timestamp 1644511149
transform 1 0 55660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2452__101
timestamp 1644511149
transform 1 0 13248 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2453__102
timestamp 1644511149
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2454__103
timestamp 1644511149
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2455__104
timestamp 1644511149
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2457_
timestamp 1644511149
transform 1 0 1932 0 -1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2458_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2459_
timestamp 1644511149
transform 1 0 1932 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2460_
timestamp 1644511149
transform 1 0 54004 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2461_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2462_
timestamp 1644511149
transform 1 0 56304 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2463_
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2464_
timestamp 1644511149
transform 1 0 56304 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2465_
timestamp 1644511149
transform 1 0 55476 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2466_
timestamp 1644511149
transform 1 0 56304 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2467_
timestamp 1644511149
transform 1 0 26680 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2468_
timestamp 1644511149
transform 1 0 56304 0 1 54400
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2469_
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2470_
timestamp 1644511149
transform 1 0 32108 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2471_
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2472_
timestamp 1644511149
transform 1 0 56304 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2473_
timestamp 1644511149
transform 1 0 56304 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2474_
timestamp 1644511149
transform 1 0 8648 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2475_
timestamp 1644511149
transform 1 0 56304 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2476_
timestamp 1644511149
transform 1 0 2208 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2477_
timestamp 1644511149
transform 1 0 56304 0 1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2478_
timestamp 1644511149
transform 1 0 35696 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2479_
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2480_
timestamp 1644511149
transform 1 0 56304 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2481_
timestamp 1644511149
transform 1 0 1932 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2482_
timestamp 1644511149
transform 1 0 56304 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2483_
timestamp 1644511149
transform 1 0 1932 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2484_
timestamp 1644511149
transform 1 0 52900 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2485_
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2486_
timestamp 1644511149
transform 1 0 56304 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2487_
timestamp 1644511149
transform 1 0 56304 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2488_
timestamp 1644511149
transform 1 0 55476 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2489_
timestamp 1644511149
transform 1 0 39652 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2490_
timestamp 1644511149
transform 1 0 8004 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2491_
timestamp 1644511149
transform 1 0 2208 0 -1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2492_
timestamp 1644511149
transform 1 0 56304 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2493_
timestamp 1644511149
transform 1 0 27968 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2494_
timestamp 1644511149
transform 1 0 56304 0 1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2495_
timestamp 1644511149
transform 1 0 1932 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2496_
timestamp 1644511149
transform 1 0 22816 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2497_
timestamp 1644511149
transform 1 0 2208 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2498_
timestamp 1644511149
transform 1 0 56304 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2499_
timestamp 1644511149
transform 1 0 1932 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2500_
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2501_
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2502_
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2503_
timestamp 1644511149
transform 1 0 8464 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2504_
timestamp 1644511149
transform 1 0 56304 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2505_
timestamp 1644511149
transform 1 0 52900 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2506_
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2507_
timestamp 1644511149
transform 1 0 24564 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2508_
timestamp 1644511149
transform 1 0 47748 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2509_
timestamp 1644511149
transform 1 0 27140 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2510_
timestamp 1644511149
transform 1 0 38272 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2511_
timestamp 1644511149
transform 1 0 56304 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2512_
timestamp 1644511149
transform 1 0 32108 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2513_
timestamp 1644511149
transform 1 0 42596 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2514_
timestamp 1644511149
transform 1 0 1932 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2515_
timestamp 1644511149
transform 1 0 46184 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2516_
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2517_
timestamp 1644511149
transform 1 0 56304 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2518_
timestamp 1644511149
transform 1 0 1932 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2519_
timestamp 1644511149
transform 1 0 1932 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2520_
timestamp 1644511149
transform 1 0 2300 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2521_
timestamp 1644511149
transform 1 0 56304 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2522_
timestamp 1644511149
transform 1 0 56304 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2523_
timestamp 1644511149
transform 1 0 56304 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2524_
timestamp 1644511149
transform 1 0 19044 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2525_
timestamp 1644511149
transform 1 0 56304 0 1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2526_
timestamp 1644511149
transform 1 0 29808 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2527_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2528_
timestamp 1644511149
transform 1 0 49496 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2529_
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2530_
timestamp 1644511149
transform 1 0 56304 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2531_
timestamp 1644511149
transform 1 0 2208 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2532_
timestamp 1644511149
transform 1 0 56304 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2533_
timestamp 1644511149
transform 1 0 15732 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2534_
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2535_
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2536_
timestamp 1644511149
transform 1 0 1932 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2537_
timestamp 1644511149
transform 1 0 56304 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2538_
timestamp 1644511149
transform 1 0 56304 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2539_
timestamp 1644511149
transform 1 0 56304 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2540_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2541_
timestamp 1644511149
transform 1 0 16744 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2542_
timestamp 1644511149
transform 1 0 55476 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2543_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2544_
timestamp 1644511149
transform 1 0 42412 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2545_
timestamp 1644511149
transform 1 0 17664 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2546_
timestamp 1644511149
transform 1 0 56304 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2547_
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2548_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2549_
timestamp 1644511149
transform 1 0 29992 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2550_
timestamp 1644511149
transform 1 0 31280 0 1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2551_
timestamp 1644511149
transform 1 0 55476 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2552_
timestamp 1644511149
transform 1 0 56304 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2553_
timestamp 1644511149
transform 1 0 35604 0 1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2554_
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2555_
timestamp 1644511149
transform 1 0 56304 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2556_
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2557_
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2558_
timestamp 1644511149
transform 1 0 1932 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2559_
timestamp 1644511149
transform 1 0 55476 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2560_
timestamp 1644511149
transform 1 0 13248 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2561_
timestamp 1644511149
transform 1 0 1932 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2562_
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2563_
timestamp 1644511149
transform 1 0 1932 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 28244 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 25760 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 29624 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 27140 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26404 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 32476 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 32752 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 24840 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 30452 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 33580 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 57868 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 10396 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  input6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 57224 0 1 9792
box -38 -48 1050 592
<< labels >>
rlabel metal3 s 0 55708 800 55948 6 active
port 0 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 33478 59200 33590 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 634 59200 746 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 59200 50268 60000 50508 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 22530 59200 22642 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 59200 52308 60000 52548 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 59200 4708 60000 4948 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 12870 59200 12982 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 14802 59200 14914 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 51510 0 51622 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 59200 18308 60000 18548 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 11582 59200 11694 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 8362 59200 8474 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 45070 0 45182 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 59200 12868 60000 13108 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 59882 59200 59994 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 59200 23068 60000 23308 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 52988 800 53228 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 45714 59200 45826 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 52154 59200 52266 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 59200 37348 60000 37588 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 53442 59200 53554 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 34766 59200 34878 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 59200 35988 60000 36228 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 59200 57068 60000 57308 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 59200 39388 60000 39628 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 10294 59200 10406 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 io_oeb[0]
port 39 nsew signal bidirectional
rlabel metal3 s 0 20348 800 20588 6 io_oeb[10]
port 40 nsew signal bidirectional
rlabel metal3 s 59200 33948 60000 34188 6 io_oeb[11]
port 41 nsew signal bidirectional
rlabel metal3 s 59200 17628 60000 17868 6 io_oeb[12]
port 42 nsew signal bidirectional
rlabel metal3 s 59200 16268 60000 16508 6 io_oeb[13]
port 43 nsew signal bidirectional
rlabel metal3 s 0 5388 800 5628 6 io_oeb[14]
port 44 nsew signal bidirectional
rlabel metal2 s 17378 59200 17490 60000 6 io_oeb[15]
port 45 nsew signal bidirectional
rlabel metal3 s 59200 1988 60000 2228 6 io_oeb[16]
port 46 nsew signal bidirectional
rlabel metal2 s 16090 0 16202 800 6 io_oeb[17]
port 47 nsew signal bidirectional
rlabel metal2 s 43782 59200 43894 60000 6 io_oeb[18]
port 48 nsew signal bidirectional
rlabel metal2 s 18022 59200 18134 60000 6 io_oeb[19]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 0 47114 800 6 io_oeb[1]
port 50 nsew signal bidirectional
rlabel metal3 s 59200 25788 60000 26028 6 io_oeb[20]
port 51 nsew signal bidirectional
rlabel metal2 s 2566 59200 2678 60000 6 io_oeb[21]
port 52 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 io_oeb[22]
port 53 nsew signal bidirectional
rlabel metal2 s 30258 59200 30370 60000 6 io_oeb[23]
port 54 nsew signal bidirectional
rlabel metal2 s 31546 59200 31658 60000 6 io_oeb[24]
port 55 nsew signal bidirectional
rlabel metal2 s 57306 0 57418 800 6 io_oeb[25]
port 56 nsew signal bidirectional
rlabel metal3 s 59200 46868 60000 47108 6 io_oeb[26]
port 57 nsew signal bidirectional
rlabel metal2 s 36054 59200 36166 60000 6 io_oeb[27]
port 58 nsew signal bidirectional
rlabel metal2 s 50222 0 50334 800 6 io_oeb[28]
port 59 nsew signal bidirectional
rlabel metal3 s 59200 38708 60000 38948 6 io_oeb[29]
port 60 nsew signal bidirectional
rlabel metal2 s 50222 59200 50334 60000 6 io_oeb[2]
port 61 nsew signal bidirectional
rlabel metal2 s 3854 59200 3966 60000 6 io_oeb[30]
port 62 nsew signal bidirectional
rlabel metal2 s 49578 0 49690 800 6 io_oeb[31]
port 63 nsew signal bidirectional
rlabel metal3 s 0 29868 800 30108 6 io_oeb[32]
port 64 nsew signal bidirectional
rlabel metal2 s 58594 0 58706 800 6 io_oeb[33]
port 65 nsew signal bidirectional
rlabel metal2 s 13514 59200 13626 60000 6 io_oeb[34]
port 66 nsew signal bidirectional
rlabel metal3 s 0 26468 800 26708 6 io_oeb[35]
port 67 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 io_oeb[36]
port 68 nsew signal bidirectional
rlabel metal3 s 0 21708 800 21948 6 io_oeb[37]
port 69 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 io_oeb[3]
port 70 nsew signal bidirectional
rlabel metal3 s 59200 -52 60000 188 6 io_oeb[4]
port 71 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 io_oeb[5]
port 72 nsew signal bidirectional
rlabel metal3 s 59200 21028 60000 21268 6 io_oeb[6]
port 73 nsew signal bidirectional
rlabel metal2 s 16090 59200 16202 60000 6 io_oeb[7]
port 74 nsew signal bidirectional
rlabel metal2 s 5142 0 5254 800 6 io_oeb[8]
port 75 nsew signal bidirectional
rlabel metal2 s 12870 0 12982 800 6 io_oeb[9]
port 76 nsew signal bidirectional
rlabel metal3 s 59200 55708 60000 55948 6 io_out[0]
port 77 nsew signal bidirectional
rlabel metal3 s 59200 32588 60000 32828 6 io_out[10]
port 78 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 io_out[11]
port 79 nsew signal bidirectional
rlabel metal3 s 0 8788 800 9028 6 io_out[12]
port 80 nsew signal bidirectional
rlabel metal2 s 48290 0 48402 800 6 io_out[13]
port 81 nsew signal bidirectional
rlabel metal3 s 59200 47548 60000 47788 6 io_out[14]
port 82 nsew signal bidirectional
rlabel metal3 s 0 49588 800 49828 6 io_out[15]
port 83 nsew signal bidirectional
rlabel metal3 s 59200 31228 60000 31468 6 io_out[16]
port 84 nsew signal bidirectional
rlabel metal2 s 56018 59200 56130 60000 6 io_out[17]
port 85 nsew signal bidirectional
rlabel metal2 s 56018 0 56130 800 6 io_out[18]
port 86 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 io_out[19]
port 87 nsew signal bidirectional
rlabel metal2 s 40562 59200 40674 60000 6 io_out[1]
port 88 nsew signal bidirectional
rlabel metal2 s 48934 59200 49046 60000 6 io_out[20]
port 89 nsew signal bidirectional
rlabel metal3 s 0 48908 800 49148 6 io_out[21]
port 90 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 io_out[22]
port 91 nsew signal bidirectional
rlabel metal3 s 59200 26468 60000 26708 6 io_out[23]
port 92 nsew signal bidirectional
rlabel metal2 s 32834 0 32946 800 6 io_out[24]
port 93 nsew signal bidirectional
rlabel metal2 s 44426 59200 44538 60000 6 io_out[25]
port 94 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 io_out[26]
port 95 nsew signal bidirectional
rlabel metal2 s 47002 59200 47114 60000 6 io_out[27]
port 96 nsew signal bidirectional
rlabel metal2 s 20598 0 20710 800 6 io_out[28]
port 97 nsew signal bidirectional
rlabel metal3 s 59200 1308 60000 1548 6 io_out[29]
port 98 nsew signal bidirectional
rlabel metal2 s 8362 0 8474 800 6 io_out[2]
port 99 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 io_out[30]
port 100 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 io_out[31]
port 101 nsew signal bidirectional
rlabel metal3 s 0 57068 800 57308 6 io_out[32]
port 102 nsew signal bidirectional
rlabel metal3 s 59200 8108 60000 8348 6 io_out[33]
port 103 nsew signal bidirectional
rlabel metal3 s 59200 48908 60000 49148 6 io_out[34]
port 104 nsew signal bidirectional
rlabel metal3 s 59200 45508 60000 45748 6 io_out[35]
port 105 nsew signal bidirectional
rlabel metal2 s 19310 59200 19422 60000 6 io_out[36]
port 106 nsew signal bidirectional
rlabel metal3 s 59200 53668 60000 53908 6 io_out[37]
port 107 nsew signal bidirectional
rlabel metal3 s 0 52308 800 52548 6 io_out[3]
port 108 nsew signal bidirectional
rlabel metal3 s 59200 34628 60000 34868 6 io_out[4]
port 109 nsew signal bidirectional
rlabel metal2 s 28326 59200 28438 60000 6 io_out[5]
port 110 nsew signal bidirectional
rlabel metal2 s 57950 59200 58062 60000 6 io_out[6]
port 111 nsew signal bidirectional
rlabel metal3 s 0 24428 800 24668 6 io_out[7]
port 112 nsew signal bidirectional
rlabel metal2 s 23174 0 23286 800 6 io_out[8]
port 113 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 io_out[9]
port 114 nsew signal bidirectional
rlabel metal3 s 59200 9468 60000 9708 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 59200 6748 60000 6988 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 20598 59200 20710 60000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 37986 59200 38098 60000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 28970 59200 29082 60000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 52798 0 52910 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 21242 59200 21354 60000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 44148 800 44388 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 59238 59200 59350 60000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 59200 10148 60000 10388 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 46188 800 46428 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 59200 3348 60000 3588 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal2 s 1278 59200 1390 60000 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 51510 59200 51622 60000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 59200 29188 60000 29428 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 23818 59200 23930 60000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 25106 59200 25218 60000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 41428 800 41668 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la1_data_out[0]
port 147 nsew signal bidirectional
rlabel metal3 s 59200 14228 60000 14468 6 la1_data_out[10]
port 148 nsew signal bidirectional
rlabel metal2 s 27038 0 27150 800 6 la1_data_out[11]
port 149 nsew signal bidirectional
rlabel metal3 s 59200 55028 60000 55268 6 la1_data_out[12]
port 150 nsew signal bidirectional
rlabel metal2 s 5786 59200 5898 60000 6 la1_data_out[13]
port 151 nsew signal bidirectional
rlabel metal2 s 32834 59200 32946 60000 6 la1_data_out[14]
port 152 nsew signal bidirectional
rlabel metal3 s 0 1988 800 2228 6 la1_data_out[15]
port 153 nsew signal bidirectional
rlabel metal3 s 59200 19668 60000 19908 6 la1_data_out[16]
port 154 nsew signal bidirectional
rlabel metal3 s 59200 42788 60000 43028 6 la1_data_out[17]
port 155 nsew signal bidirectional
rlabel metal2 s 7074 59200 7186 60000 6 la1_data_out[18]
port 156 nsew signal bidirectional
rlabel metal3 s 59200 30548 60000 30788 6 la1_data_out[19]
port 157 nsew signal bidirectional
rlabel metal3 s 0 54348 800 54588 6 la1_data_out[1]
port 158 nsew signal bidirectional
rlabel metal3 s 0 12188 800 12428 6 la1_data_out[20]
port 159 nsew signal bidirectional
rlabel metal3 s 59200 50948 60000 51188 6 la1_data_out[21]
port 160 nsew signal bidirectional
rlabel metal2 s 36698 59200 36810 60000 6 la1_data_out[22]
port 161 nsew signal bidirectional
rlabel metal2 s 15446 0 15558 800 6 la1_data_out[23]
port 162 nsew signal bidirectional
rlabel metal3 s 59200 22388 60000 22628 6 la1_data_out[24]
port 163 nsew signal bidirectional
rlabel metal3 s 0 4028 800 4268 6 la1_data_out[25]
port 164 nsew signal bidirectional
rlabel metal3 s 59200 6068 60000 6308 6 la1_data_out[26]
port 165 nsew signal bidirectional
rlabel metal3 s 0 57748 800 57988 6 la1_data_out[27]
port 166 nsew signal bidirectional
rlabel metal2 s 54086 0 54198 800 6 la1_data_out[28]
port 167 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[29]
port 168 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la1_data_out[2]
port 169 nsew signal bidirectional
rlabel metal3 s 59200 14908 60000 15148 6 la1_data_out[30]
port 170 nsew signal bidirectional
rlabel metal3 s 59200 58428 60000 58668 6 la1_data_out[31]
port 171 nsew signal bidirectional
rlabel metal3 s 0 11508 800 11748 6 la1_data_out[3]
port 172 nsew signal bidirectional
rlabel metal2 s 54730 0 54842 800 6 la1_data_out[4]
port 173 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 174 nsew signal bidirectional
rlabel metal3 s 59200 24428 60000 24668 6 la1_data_out[6]
port 175 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal bidirectional
rlabel metal3 s 59200 44148 60000 44388 6 la1_data_out[8]
port 177 nsew signal bidirectional
rlabel metal2 s 56662 59200 56774 60000 6 la1_data_out[9]
port 178 nsew signal bidirectional
rlabel metal2 s 59238 0 59350 800 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 54730 59200 54842 60000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s 5142 59200 5254 60000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 27038 59200 27150 60000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 39274 59200 39386 60000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 25750 59200 25862 60000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 48290 59200 48402 60000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 59200 11508 60000 11748 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 59200 42108 60000 42348 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 59200 40748 60000 40988 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 42494 59200 42606 60000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 41206 59200 41318 60000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 59108 800 59348 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 9650 59200 9762 60000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 41850 0 41962 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 50948 800 51188 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 211 nsew power input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 211 nsew power input
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 212 nsew ground input
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 212 nsew ground input
rlabel metal3 s 59200 27828 60000 28068 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
